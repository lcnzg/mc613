library ieee;
use ieee.std_logic_1164.all;

entity sine_wave is
	port (
		indice: in integer range 0 to 7999;
		amplitude: out integer range -2097152 to 2097152
);
end sine_wave;

architecture rtl of sine_wave is

begin

	-- lookup table
	with indice select
			amplitude <=	0 when 0,
	1647 when 1,
	3294 when 2,
	4941 when 3,
	6588 when 4,
	8235 when 5,
	9883 when 6,
	11530 when 7,
	13177 when 8,
	14824 when 9,
	16471 when 10,
	18118 when 11,
	19765 when 12,
	21412 when 13,
	23059 when 14,
	24706 when 15,
	26353 when 16,
	28000 when 17,
	29647 when 18,
	31294 when 19,
	32941 when 20,
	34588 when 21,
	36234 when 22,
	37881 when 23,
	39528 when 24,
	41175 when 25,
	42822 when 26,
	44468 when 27,
	46115 when 28,
	47762 when 29,
	49408 when 30,
	51055 when 31,
	52702 when 32,
	54348 when 33,
	55995 when 34,
	57641 when 35,
	59288 when 36,
	60934 when 37,
	62580 when 38,
	64227 when 39,
	65873 when 40,
	67519 when 41,
	69166 when 42,
	70812 when 43,
	72458 when 44,
	74104 when 45,
	75750 when 46,
	77396 when 47,
	79042 when 48,
	80688 when 49,
	82334 when 50,
	83980 when 51,
	85625 when 52,
	87271 when 53,
	88917 when 54,
	90562 when 55,
	92208 when 56,
	93853 when 57,
	95499 when 58,
	97144 when 59,
	98789 when 60,
	100435 when 61,
	102080 when 62,
	103725 when 63,
	105370 when 64,
	107015 when 65,
	108660 when 66,
	110305 when 67,
	111950 when 68,
	113594 when 69,
	115239 when 70,
	116883 when 71,
	118528 when 72,
	120172 when 73,
	121817 when 74,
	123461 when 75,
	125105 when 76,
	126749 when 77,
	128393 when 78,
	130037 when 79,
	131681 when 80,
	133325 when 81,
	134969 when 82,
	136612 when 83,
	138256 when 84,
	139899 when 85,
	141543 when 86,
	143186 when 87,
	144829 when 88,
	146472 when 89,
	148116 when 90,
	149758 when 91,
	151401 when 92,
	153044 when 93,
	154687 when 94,
	156329 when 95,
	157972 when 96,
	159614 when 97,
	161256 when 98,
	162899 when 99,
	164541 when 100,
	166183 when 101,
	167824 when 102,
	169466 when 103,
	171108 when 104,
	172749 when 105,
	174391 when 106,
	176032 when 107,
	177673 when 108,
	179315 when 109,
	180956 when 110,
	182597 when 111,
	184237 when 112,
	185878 when 113,
	187519 when 114,
	189159 when 115,
	190799 when 116,
	192440 when 117,
	194080 when 118,
	195720 when 119,
	197359 when 120,
	198999 when 121,
	200639 when 122,
	202278 when 123,
	203918 when 124,
	205557 when 125,
	207196 when 126,
	208835 when 127,
	210474 when 128,
	212112 when 129,
	213751 when 130,
	215390 when 131,
	217028 when 132,
	218666 when 133,
	220304 when 134,
	221942 when 135,
	223580 when 136,
	225217 when 137,
	226855 when 138,
	228492 when 139,
	230130 when 140,
	231767 when 141,
	233404 when 142,
	235040 when 143,
	236677 when 144,
	238313 when 145,
	239950 when 146,
	241586 when 147,
	243222 when 148,
	244858 when 149,
	246494 when 150,
	248129 when 151,
	249765 when 152,
	251400 when 153,
	253035 when 154,
	254670 when 155,
	256305 when 156,
	257940 when 157,
	259574 when 158,
	261209 when 159,
	262843 when 160,
	264477 when 161,
	266111 when 162,
	267744 when 163,
	269378 when 164,
	271011 when 165,
	272645 when 166,
	274278 when 167,
	275910 when 168,
	277543 when 169,
	279176 when 170,
	280808 when 171,
	282440 when 172,
	284072 when 173,
	285704 when 174,
	287336 when 175,
	288967 when 176,
	290598 when 177,
	292230 when 178,
	293861 when 179,
	295491 when 180,
	297122 when 181,
	298752 when 182,
	300382 when 183,
	302013 when 184,
	303642 when 185,
	305272 when 186,
	306901 when 187,
	308531 when 188,
	310160 when 189,
	311789 when 190,
	313417 when 191,
	315046 when 192,
	316674 when 193,
	318302 when 194,
	319930 when 195,
	321558 when 196,
	323185 when 197,
	324813 when 198,
	326440 when 199,
	328067 when 200,
	329694 when 201,
	331320 when 202,
	332946 when 203,
	334573 when 204,
	336198 when 205,
	337824 when 206,
	339450 when 207,
	341075 when 208,
	342700 when 209,
	344325 when 210,
	345949 when 211,
	347574 when 212,
	349198 when 213,
	350822 when 214,
	352446 when 215,
	354069 when 216,
	355693 when 217,
	357316 when 218,
	358939 when 219,
	360561 when 220,
	362184 when 221,
	363806 when 222,
	365428 when 223,
	367050 when 224,
	368672 when 225,
	370293 when 226,
	371914 when 227,
	373535 when 228,
	375155 when 229,
	376776 when 230,
	378396 when 231,
	380016 when 232,
	381636 when 233,
	383255 when 234,
	384874 when 235,
	386493 when 236,
	388112 when 237,
	389731 when 238,
	391349 when 239,
	392967 when 240,
	394585 when 241,
	396202 when 242,
	397820 when 243,
	399437 when 244,
	401054 when 245,
	402670 when 246,
	404287 when 247,
	405903 when 248,
	407518 when 249,
	409134 when 250,
	410749 when 251,
	412364 when 252,
	413979 when 253,
	415594 when 254,
	417208 when 255,
	418822 when 256,
	420436 when 257,
	422050 when 258,
	423663 when 259,
	425276 when 260,
	426889 when 261,
	428501 when 262,
	430113 when 263,
	431725 when 264,
	433337 when 265,
	434948 when 266,
	436559 when 267,
	438170 when 268,
	439781 when 269,
	441391 when 270,
	443001 when 271,
	444611 when 272,
	446221 when 273,
	447830 when 274,
	449439 when 275,
	451048 when 276,
	452656 when 277,
	454264 when 278,
	455872 when 279,
	457480 when 280,
	459087 when 281,
	460694 when 282,
	462301 when 283,
	463907 when 284,
	465513 when 285,
	467119 when 286,
	468725 when 287,
	470330 when 288,
	471935 when 289,
	473540 when 290,
	475144 when 291,
	476748 when 292,
	478352 when 293,
	479955 when 294,
	481559 when 295,
	483162 when 296,
	484764 when 297,
	486367 when 298,
	487969 when 299,
	489570 when 300,
	491172 when 301,
	492773 when 302,
	494374 when 303,
	495974 when 304,
	497575 when 305,
	499174 when 306,
	500774 when 307,
	502373 when 308,
	503972 when 309,
	505571 when 310,
	507169 when 311,
	508767 when 312,
	510365 when 313,
	511963 when 314,
	513560 when 315,
	515157 when 316,
	516753 when 317,
	518349 when 318,
	519945 when 319,
	521540 when 320,
	523136 when 321,
	524731 when 322,
	526325 when 323,
	527919 when 324,
	529513 when 325,
	531107 when 326,
	532700 when 327,
	534293 when 328,
	535886 when 329,
	537478 when 330,
	539070 when 331,
	540661 when 332,
	542253 when 333,
	543843 when 334,
	545434 when 335,
	547024 when 336,
	548614 when 337,
	550204 when 338,
	551793 when 339,
	553382 when 340,
	554970 when 341,
	556559 when 342,
	558147 when 343,
	559734 when 344,
	561321 when 345,
	562908 when 346,
	564495 when 347,
	566081 when 348,
	567666 when 349,
	569252 when 350,
	570837 when 351,
	572422 when 352,
	574006 when 353,
	575590 when 354,
	577174 when 355,
	578757 when 356,
	580340 when 357,
	581923 when 358,
	583505 when 359,
	585087 when 360,
	586668 when 361,
	588249 when 362,
	589830 when 363,
	591411 when 364,
	592991 when 365,
	594570 when 366,
	596150 when 367,
	597729 when 368,
	599307 when 369,
	600886 when 370,
	602463 when 371,
	604041 when 372,
	605618 when 373,
	607195 when 374,
	608771 when 375,
	610347 when 376,
	611923 when 377,
	613498 when 378,
	615073 when 379,
	616647 when 380,
	618221 when 381,
	619795 when 382,
	621368 when 383,
	622941 when 384,
	624514 when 385,
	626086 when 386,
	627658 when 387,
	629229 when 388,
	630800 when 389,
	632371 when 390,
	633941 when 391,
	635511 when 392,
	637080 when 393,
	638650 when 394,
	640218 when 395,
	641786 when 396,
	643354 when 397,
	644922 when 398,
	646489 when 399,
	648056 when 400,
	649622 when 401,
	651188 when 402,
	652753 when 403,
	654318 when 404,
	655883 when 405,
	657447 when 406,
	659011 when 407,
	660575 when 408,
	662138 when 409,
	663700 when 410,
	665263 when 411,
	666824 when 412,
	668386 when 413,
	669947 when 414,
	671507 when 415,
	673068 when 416,
	674627 when 417,
	676187 when 418,
	677746 when 419,
	679304 when 420,
	680862 when 421,
	682420 when 422,
	683977 when 423,
	685534 when 424,
	687090 when 425,
	688646 when 426,
	690202 when 427,
	691757 when 428,
	693312 when 429,
	694866 when 430,
	696420 when 431,
	697973 when 432,
	699526 when 433,
	701079 when 434,
	702631 when 435,
	704183 when 436,
	705734 when 437,
	707285 when 438,
	708835 when 439,
	710385 when 440,
	711934 when 441,
	713483 when 442,
	715032 when 443,
	716580 when 444,
	718128 when 445,
	719675 when 446,
	721222 when 447,
	722769 when 448,
	724315 when 449,
	725860 when 450,
	727405 when 451,
	728950 when 452,
	730494 when 453,
	732038 when 454,
	733581 when 455,
	735124 when 456,
	736666 when 457,
	738208 when 458,
	739749 when 459,
	741290 when 460,
	742831 when 461,
	744371 when 462,
	745911 when 463,
	747450 when 464,
	748989 when 465,
	750527 when 466,
	752065 when 467,
	753602 when 468,
	755139 when 469,
	756675 when 470,
	758211 when 471,
	759747 when 472,
	761281 when 473,
	762816 when 474,
	764350 when 475,
	765884 when 476,
	767417 when 477,
	768949 when 478,
	770481 when 479,
	772013 when 480,
	773544 when 481,
	775075 when 482,
	776605 when 483,
	778135 when 484,
	779664 when 485,
	781193 when 486,
	782721 when 487,
	784249 when 488,
	785777 when 489,
	787304 when 490,
	788830 when 491,
	790356 when 492,
	791881 when 493,
	793406 when 494,
	794931 when 495,
	796454 when 496,
	797978 when 497,
	799501 when 498,
	801023 when 499,
	802545 when 500,
	804067 when 501,
	805588 when 502,
	807108 when 503,
	808628 when 504,
	810148 when 505,
	811667 when 506,
	813185 when 507,
	814703 when 508,
	816221 when 509,
	817738 when 510,
	819254 when 511,
	820770 when 512,
	822286 when 513,
	823800 when 514,
	825315 when 515,
	826829 when 516,
	828342 when 517,
	829855 when 518,
	831368 when 519,
	832879 when 520,
	834391 when 521,
	835902 when 522,
	837412 when 523,
	838922 when 524,
	840431 when 525,
	841940 when 526,
	843448 when 527,
	844956 when 528,
	846463 when 529,
	847970 when 530,
	849476 when 531,
	850982 when 532,
	852487 when 533,
	853992 when 534,
	855496 when 535,
	856999 when 536,
	858502 when 537,
	860005 when 538,
	861507 when 539,
	863008 when 540,
	864509 when 541,
	866009 when 542,
	867509 when 543,
	869009 when 544,
	870507 when 545,
	872006 when 546,
	873503 when 547,
	875000 when 548,
	876497 when 549,
	877993 when 550,
	879489 when 551,
	880984 when 552,
	882478 when 553,
	883972 when 554,
	885465 when 555,
	886958 when 556,
	888450 when 557,
	889942 when 558,
	891433 when 559,
	892924 when 560,
	894414 when 561,
	895903 when 562,
	897392 when 563,
	898881 when 564,
	900369 when 565,
	901856 when 566,
	903343 when 567,
	904829 when 568,
	906315 when 569,
	907800 when 570,
	909284 when 571,
	910768 when 572,
	912251 when 573,
	913734 when 574,
	915217 when 575,
	916698 when 576,
	918179 when 577,
	919660 when 578,
	921140 when 579,
	922619 when 580,
	924098 when 581,
	925576 when 582,
	927054 when 583,
	928531 when 584,
	930008 when 585,
	931484 when 586,
	932959 when 587,
	934434 when 588,
	935908 when 589,
	937382 when 590,
	938855 when 591,
	940328 when 592,
	941800 when 593,
	943271 when 594,
	944742 when 595,
	946212 when 596,
	947682 when 597,
	949151 when 598,
	950619 when 599,
	952087 when 600,
	953554 when 601,
	955021 when 602,
	956487 when 603,
	957953 when 604,
	959418 when 605,
	960882 when 606,
	962346 when 607,
	963809 when 608,
	965271 when 609,
	966733 when 610,
	968195 when 611,
	969655 when 612,
	971116 when 613,
	972575 when 614,
	974034 when 615,
	975493 when 616,
	976950 when 617,
	978407 when 618,
	979864 when 619,
	981320 when 620,
	982775 when 621,
	984230 when 622,
	985684 when 623,
	987138 when 624,
	988591 when 625,
	990043 when 626,
	991495 when 627,
	992946 when 628,
	994396 when 629,
	995846 when 630,
	997295 when 631,
	998744 when 632,
	1000192 when 633,
	1001639 when 634,
	1003086 when 635,
	1004532 when 636,
	1005978 when 637,
	1007423 when 638,
	1008867 when 639,
	1010311 when 640,
	1011754 when 641,
	1013196 when 642,
	1014638 when 643,
	1016079 when 644,
	1017520 when 645,
	1018960 when 646,
	1020399 when 647,
	1021838 when 648,
	1023276 when 649,
	1024713 when 650,
	1026150 when 651,
	1027586 when 652,
	1029021 when 653,
	1030456 when 654,
	1031891 when 655,
	1033324 when 656,
	1034757 when 657,
	1036189 when 658,
	1037621 when 659,
	1039052 when 660,
	1040483 when 661,
	1041912 when 662,
	1043341 when 663,
	1044770 when 664,
	1046198 when 665,
	1047625 when 666,
	1049051 when 667,
	1050477 when 668,
	1051903 when 669,
	1053327 when 670,
	1054751 when 671,
	1056174 when 672,
	1057597 when 673,
	1059019 when 674,
	1060440 when 675,
	1061861 when 676,
	1063281 when 677,
	1064700 when 678,
	1066119 when 679,
	1067537 when 680,
	1068955 when 681,
	1070371 when 682,
	1071787 when 683,
	1073203 when 684,
	1074618 when 685,
	1076032 when 686,
	1077445 when 687,
	1078858 when 688,
	1080270 when 689,
	1081681 when 690,
	1083092 when 691,
	1084502 when 692,
	1085912 when 693,
	1087320 when 694,
	1088729 when 695,
	1090136 when 696,
	1091543 when 697,
	1092949 when 698,
	1094354 when 699,
	1095759 when 700,
	1097163 when 701,
	1098566 when 702,
	1099969 when 703,
	1101371 when 704,
	1102772 when 705,
	1104173 when 706,
	1105573 when 707,
	1106972 when 708,
	1108371 when 709,
	1109769 when 710,
	1111166 when 711,
	1112563 when 712,
	1113958 when 713,
	1115354 when 714,
	1116748 when 715,
	1118142 when 716,
	1119535 when 717,
	1120927 when 718,
	1122319 when 719,
	1123710 when 720,
	1125101 when 721,
	1126490 when 722,
	1127879 when 723,
	1129267 when 724,
	1130655 when 725,
	1132042 when 726,
	1133428 when 727,
	1134814 when 728,
	1136198 when 729,
	1137582 when 730,
	1138966 when 731,
	1140348 when 732,
	1141730 when 733,
	1143112 when 734,
	1144492 when 735,
	1145872 when 736,
	1147251 when 737,
	1148630 when 738,
	1150007 when 739,
	1151384 when 740,
	1152761 when 741,
	1154136 when 742,
	1155511 when 743,
	1156885 when 744,
	1158259 when 745,
	1159631 when 746,
	1161003 when 747,
	1162375 when 748,
	1163745 when 749,
	1165115 when 750,
	1166484 when 751,
	1167853 when 752,
	1169221 when 753,
	1170588 when 754,
	1171954 when 755,
	1173319 when 756,
	1174684 when 757,
	1176048 when 758,
	1177412 when 759,
	1178774 when 760,
	1180136 when 761,
	1181497 when 762,
	1182858 when 763,
	1184218 when 764,
	1185577 when 765,
	1186935 when 766,
	1188292 when 767,
	1189649 when 768,
	1191005 when 769,
	1192361 when 770,
	1193715 when 771,
	1195069 when 772,
	1196422 when 773,
	1197775 when 774,
	1199126 when 775,
	1200477 when 776,
	1201827 when 777,
	1203177 when 778,
	1204525 when 779,
	1205873 when 780,
	1207221 when 781,
	1208567 when 782,
	1209913 when 783,
	1211258 when 784,
	1212602 when 785,
	1213945 when 786,
	1215288 when 787,
	1216630 when 788,
	1217971 when 789,
	1219312 when 790,
	1220652 when 791,
	1221991 when 792,
	1223329 when 793,
	1224666 when 794,
	1226003 when 795,
	1227339 when 796,
	1228674 when 797,
	1230008 when 798,
	1231342 when 799,
	1232675 when 800,
	1234007 when 801,
	1235339 when 802,
	1236669 when 803,
	1237999 when 804,
	1239328 when 805,
	1240656 when 806,
	1241984 when 807,
	1243311 when 808,
	1244637 when 809,
	1245962 when 810,
	1247287 when 811,
	1248610 when 812,
	1249933 when 813,
	1251256 when 814,
	1252577 when 815,
	1253898 when 816,
	1255218 when 817,
	1256537 when 818,
	1257855 when 819,
	1259172 when 820,
	1260489 when 821,
	1261805 when 822,
	1263120 when 823,
	1264435 when 824,
	1265749 when 825,
	1267061 when 826,
	1268374 when 827,
	1269685 when 828,
	1270995 when 829,
	1272305 when 830,
	1273614 when 831,
	1274922 when 832,
	1276230 when 833,
	1277536 when 834,
	1278842 when 835,
	1280147 when 836,
	1281451 when 837,
	1282755 when 838,
	1284057 when 839,
	1285359 when 840,
	1286660 when 841,
	1287961 when 842,
	1289260 when 843,
	1290559 when 844,
	1291857 when 845,
	1293154 when 846,
	1294450 when 847,
	1295746 when 848,
	1297040 when 849,
	1298334 when 850,
	1299627 when 851,
	1300920 when 852,
	1302211 when 853,
	1303502 when 854,
	1304792 when 855,
	1306081 when 856,
	1307369 when 857,
	1308656 when 858,
	1309943 when 859,
	1311229 when 860,
	1312514 when 861,
	1313798 when 862,
	1315082 when 863,
	1316364 when 864,
	1317646 when 865,
	1318927 when 866,
	1320207 when 867,
	1321487 when 868,
	1322765 when 869,
	1324043 when 870,
	1325320 when 871,
	1326596 when 872,
	1327871 when 873,
	1329146 when 874,
	1330419 when 875,
	1331692 when 876,
	1332964 when 877,
	1334235 when 878,
	1335505 when 879,
	1336775 when 880,
	1338044 when 881,
	1339312 when 882,
	1340579 when 883,
	1341845 when 884,
	1343110 when 885,
	1344375 when 886,
	1345639 when 887,
	1346901 when 888,
	1348164 when 889,
	1349425 when 890,
	1350685 when 891,
	1351945 when 892,
	1353203 when 893,
	1354461 when 894,
	1355718 when 895,
	1356975 when 896,
	1358230 when 897,
	1359485 when 898,
	1360738 when 899,
	1361991 when 900,
	1363243 when 901,
	1364495 when 902,
	1365745 when 903,
	1366994 when 904,
	1368243 when 905,
	1369491 when 906,
	1370738 when 907,
	1371984 when 908,
	1373229 when 909,
	1374474 when 910,
	1375717 when 911,
	1376960 when 912,
	1378202 when 913,
	1379443 when 914,
	1380683 when 915,
	1381923 when 916,
	1383161 when 917,
	1384399 when 918,
	1385636 when 919,
	1386872 when 920,
	1388107 when 921,
	1389341 when 922,
	1390574 when 923,
	1391807 when 924,
	1393038 when 925,
	1394269 when 926,
	1395499 when 927,
	1396728 when 928,
	1397956 when 929,
	1399184 when 930,
	1400410 when 931,
	1401636 when 932,
	1402861 when 933,
	1404084 when 934,
	1405307 when 935,
	1406530 when 936,
	1407751 when 937,
	1408971 when 938,
	1410191 when 939,
	1411410 when 940,
	1412627 when 941,
	1413844 when 942,
	1415060 when 943,
	1416276 when 944,
	1417490 when 945,
	1418703 when 946,
	1419916 when 947,
	1421128 when 948,
	1422338 when 949,
	1423548 when 950,
	1424757 when 951,
	1425966 when 952,
	1427173 when 953,
	1428379 when 954,
	1429585 when 955,
	1430790 when 956,
	1431993 when 957,
	1433196 when 958,
	1434398 when 959,
	1435599 when 960,
	1436800 when 961,
	1437999 when 962,
	1439197 when 963,
	1440395 when 964,
	1441592 when 965,
	1442787 when 966,
	1443982 when 967,
	1445176 when 968,
	1446370 when 969,
	1447562 when 970,
	1448753 when 971,
	1449944 when 972,
	1451133 when 973,
	1452322 when 974,
	1453510 when 975,
	1454696 when 976,
	1455882 when 977,
	1457067 when 978,
	1458252 when 979,
	1459435 when 980,
	1460617 when 981,
	1461799 when 982,
	1462979 when 983,
	1464159 when 984,
	1465338 when 985,
	1466516 when 986,
	1467693 when 987,
	1468869 when 988,
	1470044 when 989,
	1471218 when 990,
	1472391 when 991,
	1473564 when 992,
	1474735 when 993,
	1475906 when 994,
	1477076 when 995,
	1478244 when 996,
	1479412 when 997,
	1480579 when 998,
	1481745 when 999,
	1482910 when 1000,
	1484075 when 1001,
	1485238 when 1002,
	1486400 when 1003,
	1487562 when 1004,
	1488722 when 1005,
	1489882 when 1006,
	1491041 when 1007,
	1492198 when 1008,
	1493355 when 1009,
	1494511 when 1010,
	1495666 when 1011,
	1496820 when 1012,
	1497974 when 1013,
	1499126 when 1014,
	1500277 when 1015,
	1501428 when 1016,
	1502577 when 1017,
	1503726 when 1018,
	1504873 when 1019,
	1506020 when 1020,
	1507166 when 1021,
	1508311 when 1022,
	1509455 when 1023,
	1510598 when 1024,
	1511740 when 1025,
	1512881 when 1026,
	1514021 when 1027,
	1515160 when 1028,
	1516298 when 1029,
	1517436 when 1030,
	1518572 when 1031,
	1519708 when 1032,
	1520842 when 1033,
	1521976 when 1034,
	1523109 when 1035,
	1524240 when 1036,
	1525371 when 1037,
	1526501 when 1038,
	1527630 when 1039,
	1528758 when 1040,
	1529885 when 1041,
	1531011 when 1042,
	1532136 when 1043,
	1533261 when 1044,
	1534384 when 1045,
	1535506 when 1046,
	1536627 when 1047,
	1537748 when 1048,
	1538867 when 1049,
	1539986 when 1050,
	1541103 when 1051,
	1542220 when 1052,
	1543336 when 1053,
	1544451 when 1054,
	1545564 when 1055,
	1546677 when 1056,
	1547789 when 1057,
	1548900 when 1058,
	1550010 when 1059,
	1551119 when 1060,
	1552227 when 1061,
	1553334 when 1062,
	1554440 when 1063,
	1555545 when 1064,
	1556649 when 1065,
	1557753 when 1066,
	1558855 when 1067,
	1559956 when 1068,
	1561057 when 1069,
	1562156 when 1070,
	1563254 when 1071,
	1564352 when 1072,
	1565448 when 1073,
	1566544 when 1074,
	1567639 when 1075,
	1568732 when 1076,
	1569825 when 1077,
	1570916 when 1078,
	1572007 when 1079,
	1573097 when 1080,
	1574186 when 1081,
	1575273 when 1082,
	1576360 when 1083,
	1577446 when 1084,
	1578531 when 1085,
	1579615 when 1086,
	1580698 when 1087,
	1581780 when 1088,
	1582861 when 1089,
	1583941 when 1090,
	1585020 when 1091,
	1586098 when 1092,
	1587175 when 1093,
	1588251 when 1094,
	1589326 when 1095,
	1590400 when 1096,
	1591473 when 1097,
	1592546 when 1098,
	1593617 when 1099,
	1594687 when 1100,
	1595756 when 1101,
	1596824 when 1102,
	1597892 when 1103,
	1598958 when 1104,
	1600023 when 1105,
	1601087 when 1106,
	1602151 when 1107,
	1603213 when 1108,
	1604274 when 1109,
	1605335 when 1110,
	1606394 when 1111,
	1607452 when 1112,
	1608510 when 1113,
	1609566 when 1114,
	1610621 when 1115,
	1611676 when 1116,
	1612729 when 1117,
	1613782 when 1118,
	1614833 when 1119,
	1615883 when 1120,
	1616933 when 1121,
	1617981 when 1122,
	1619029 when 1123,
	1620075 when 1124,
	1621120 when 1125,
	1622165 when 1126,
	1623208 when 1127,
	1624251 when 1128,
	1625292 when 1129,
	1626332 when 1130,
	1627372 when 1131,
	1628410 when 1132,
	1629448 when 1133,
	1630484 when 1134,
	1631519 when 1135,
	1632554 when 1136,
	1633587 when 1137,
	1634619 when 1138,
	1635651 when 1139,
	1636681 when 1140,
	1637711 when 1141,
	1638739 when 1142,
	1639766 when 1143,
	1640792 when 1144,
	1641818 when 1145,
	1642842 when 1146,
	1643865 when 1147,
	1644888 when 1148,
	1645909 when 1149,
	1646929 when 1150,
	1647948 when 1151,
	1648966 when 1152,
	1649984 when 1153,
	1651000 when 1154,
	1652015 when 1155,
	1653029 when 1156,
	1654042 when 1157,
	1655054 when 1158,
	1656065 when 1159,
	1657075 when 1160,
	1658084 when 1161,
	1659092 when 1162,
	1660099 when 1163,
	1661105 when 1164,
	1662110 when 1165,
	1663114 when 1166,
	1664117 when 1167,
	1665119 when 1168,
	1666119 when 1169,
	1667119 when 1170,
	1668118 when 1171,
	1669116 when 1172,
	1670112 when 1173,
	1671108 when 1174,
	1672103 when 1175,
	1673096 when 1176,
	1674089 when 1177,
	1675080 when 1178,
	1676071 when 1179,
	1677060 when 1180,
	1678049 when 1181,
	1679036 when 1182,
	1680022 when 1183,
	1681008 when 1184,
	1681992 when 1185,
	1682975 when 1186,
	1683958 when 1187,
	1684939 when 1188,
	1685919 when 1189,
	1686898 when 1190,
	1687876 when 1191,
	1688853 when 1192,
	1689829 when 1193,
	1690804 when 1194,
	1691778 when 1195,
	1692751 when 1196,
	1693722 when 1197,
	1694693 when 1198,
	1695663 when 1199,
	1696632 when 1200,
	1697599 when 1201,
	1698566 when 1202,
	1699531 when 1203,
	1700496 when 1204,
	1701459 when 1205,
	1702422 when 1206,
	1703383 when 1207,
	1704343 when 1208,
	1705302 when 1209,
	1706261 when 1210,
	1707218 when 1211,
	1708174 when 1212,
	1709129 when 1213,
	1710083 when 1214,
	1711036 when 1215,
	1711987 when 1216,
	1712938 when 1217,
	1713888 when 1218,
	1714837 when 1219,
	1715784 when 1220,
	1716731 when 1221,
	1717676 when 1222,
	1718621 when 1223,
	1719564 when 1224,
	1720507 when 1225,
	1721448 when 1226,
	1722388 when 1227,
	1723327 when 1228,
	1724265 when 1229,
	1725202 when 1230,
	1726138 when 1231,
	1727073 when 1232,
	1728007 when 1233,
	1728940 when 1234,
	1729871 when 1235,
	1730802 when 1236,
	1731731 when 1237,
	1732660 when 1238,
	1733587 when 1239,
	1734514 when 1240,
	1735439 when 1241,
	1736363 when 1242,
	1737286 when 1243,
	1738208 when 1244,
	1739129 when 1245,
	1740049 when 1246,
	1740968 when 1247,
	1741886 when 1248,
	1742803 when 1249,
	1743718 when 1250,
	1744633 when 1251,
	1745546 when 1252,
	1746459 when 1253,
	1747370 when 1254,
	1748280 when 1255,
	1749189 when 1256,
	1750097 when 1257,
	1751004 when 1258,
	1751910 when 1259,
	1752815 when 1260,
	1753719 when 1261,
	1754622 when 1262,
	1755523 when 1263,
	1756424 when 1264,
	1757323 when 1265,
	1758221 when 1266,
	1759119 when 1267,
	1760015 when 1268,
	1760910 when 1269,
	1761804 when 1270,
	1762697 when 1271,
	1763589 when 1272,
	1764479 when 1273,
	1765369 when 1274,
	1766258 when 1275,
	1767145 when 1276,
	1768031 when 1277,
	1768917 when 1278,
	1769801 when 1279,
	1770684 when 1280,
	1771566 when 1281,
	1772447 when 1282,
	1773327 when 1283,
	1774205 when 1284,
	1775083 when 1285,
	1775960 when 1286,
	1776835 when 1287,
	1777709 when 1288,
	1778583 when 1289,
	1779455 when 1290,
	1780326 when 1291,
	1781196 when 1292,
	1782065 when 1293,
	1782933 when 1294,
	1783799 when 1295,
	1784665 when 1296,
	1785529 when 1297,
	1786393 when 1298,
	1787255 when 1299,
	1788116 when 1300,
	1788976 when 1301,
	1789835 when 1302,
	1790693 when 1303,
	1791550 when 1304,
	1792405 when 1305,
	1793260 when 1306,
	1794113 when 1307,
	1794966 when 1308,
	1795817 when 1309,
	1796667 when 1310,
	1797516 when 1311,
	1798364 when 1312,
	1799211 when 1313,
	1800056 when 1314,
	1800901 when 1315,
	1801744 when 1316,
	1802587 when 1317,
	1803428 when 1318,
	1804268 when 1319,
	1805107 when 1320,
	1805945 when 1321,
	1806782 when 1322,
	1807617 when 1323,
	1808452 when 1324,
	1809285 when 1325,
	1810117 when 1326,
	1810949 when 1327,
	1811779 when 1328,
	1812608 when 1329,
	1813436 when 1330,
	1814262 when 1331,
	1815088 when 1332,
	1815912 when 1333,
	1816736 when 1334,
	1817558 when 1335,
	1818379 when 1336,
	1819199 when 1337,
	1820018 when 1338,
	1820836 when 1339,
	1821652 when 1340,
	1822468 when 1341,
	1823282 when 1342,
	1824095 when 1343,
	1824908 when 1344,
	1825719 when 1345,
	1826528 when 1346,
	1827337 when 1347,
	1828145 when 1348,
	1828951 when 1349,
	1829757 when 1350,
	1830561 when 1351,
	1831364 when 1352,
	1832166 when 1353,
	1832967 when 1354,
	1833767 when 1355,
	1834565 when 1356,
	1835363 when 1357,
	1836159 when 1358,
	1836954 when 1359,
	1837748 when 1360,
	1838541 when 1361,
	1839333 when 1362,
	1840124 when 1363,
	1840913 when 1364,
	1841702 when 1365,
	1842489 when 1366,
	1843275 when 1367,
	1844060 when 1368,
	1844844 when 1369,
	1845627 when 1370,
	1846408 when 1371,
	1847188 when 1372,
	1847968 when 1373,
	1848746 when 1374,
	1849523 when 1375,
	1850299 when 1376,
	1851074 when 1377,
	1851847 when 1378,
	1852620 when 1379,
	1853391 when 1380,
	1854161 when 1381,
	1854930 when 1382,
	1855698 when 1383,
	1856465 when 1384,
	1857230 when 1385,
	1857995 when 1386,
	1858758 when 1387,
	1859520 when 1388,
	1860281 when 1389,
	1861041 when 1390,
	1861800 when 1391,
	1862557 when 1392,
	1863314 when 1393,
	1864069 when 1394,
	1864823 when 1395,
	1865576 when 1396,
	1866328 when 1397,
	1867078 when 1398,
	1867828 when 1399,
	1868576 when 1400,
	1869323 when 1401,
	1870069 when 1402,
	1870814 when 1403,
	1871558 when 1404,
	1872301 when 1405,
	1873042 when 1406,
	1873782 when 1407,
	1874521 when 1408,
	1875259 when 1409,
	1875996 when 1410,
	1876732 when 1411,
	1877466 when 1412,
	1878200 when 1413,
	1878932 when 1414,
	1879663 when 1415,
	1880393 when 1416,
	1881121 when 1417,
	1881849 when 1418,
	1882575 when 1419,
	1883300 when 1420,
	1884024 when 1421,
	1884747 when 1422,
	1885469 when 1423,
	1886190 when 1424,
	1886909 when 1425,
	1887627 when 1426,
	1888344 when 1427,
	1889060 when 1428,
	1889775 when 1429,
	1890488 when 1430,
	1891201 when 1431,
	1891912 when 1432,
	1892622 when 1433,
	1893331 when 1434,
	1894039 when 1435,
	1894745 when 1436,
	1895451 when 1437,
	1896155 when 1438,
	1896858 when 1439,
	1897560 when 1440,
	1898261 when 1441,
	1898960 when 1442,
	1899658 when 1443,
	1900356 when 1444,
	1901052 when 1445,
	1901747 when 1446,
	1902440 when 1447,
	1903133 when 1448,
	1903824 when 1449,
	1904514 when 1450,
	1905203 when 1451,
	1905891 when 1452,
	1906578 when 1453,
	1907263 when 1454,
	1907947 when 1455,
	1908631 when 1456,
	1909312 when 1457,
	1909993 when 1458,
	1910673 when 1459,
	1911351 when 1460,
	1912028 when 1461,
	1912704 when 1462,
	1913379 when 1463,
	1914053 when 1464,
	1914725 when 1465,
	1915397 when 1466,
	1916067 when 1467,
	1916736 when 1468,
	1917404 when 1469,
	1918070 when 1470,
	1918736 when 1471,
	1919400 when 1472,
	1920063 when 1473,
	1920725 when 1474,
	1921385 when 1475,
	1922045 when 1476,
	1922703 when 1477,
	1923360 when 1478,
	1924016 when 1479,
	1924671 when 1480,
	1925324 when 1481,
	1925977 when 1482,
	1926628 when 1483,
	1927278 when 1484,
	1927927 when 1485,
	1928574 when 1486,
	1929221 when 1487,
	1929866 when 1488,
	1930510 when 1489,
	1931153 when 1490,
	1931795 when 1491,
	1932435 when 1492,
	1933074 when 1493,
	1933712 when 1494,
	1934349 when 1495,
	1934985 when 1496,
	1935619 when 1497,
	1936253 when 1498,
	1936885 when 1499,
	1937516 when 1500,
	1938146 when 1501,
	1938774 when 1502,
	1939401 when 1503,
	1940028 when 1504,
	1940652 when 1505,
	1941276 when 1506,
	1941899 when 1507,
	1942520 when 1508,
	1943140 when 1509,
	1943759 when 1510,
	1944377 when 1511,
	1944993 when 1512,
	1945609 when 1513,
	1946223 when 1514,
	1946836 when 1515,
	1947448 when 1516,
	1948058 when 1517,
	1948668 when 1518,
	1949276 when 1519,
	1949883 when 1520,
	1950488 when 1521,
	1951093 when 1522,
	1951696 when 1523,
	1952298 when 1524,
	1952899 when 1525,
	1953499 when 1526,
	1954097 when 1527,
	1954695 when 1528,
	1955291 when 1529,
	1955886 when 1530,
	1956479 when 1531,
	1957072 when 1532,
	1957663 when 1533,
	1958253 when 1534,
	1958842 when 1535,
	1959430 when 1536,
	1960016 when 1537,
	1960601 when 1538,
	1961186 when 1539,
	1961768 when 1540,
	1962350 when 1541,
	1962930 when 1542,
	1963509 when 1543,
	1964087 when 1544,
	1964664 when 1545,
	1965240 when 1546,
	1965814 when 1547,
	1966387 when 1548,
	1966959 when 1549,
	1967530 when 1550,
	1968099 when 1551,
	1968668 when 1552,
	1969235 when 1553,
	1969800 when 1554,
	1970365 when 1555,
	1970929 when 1556,
	1971491 when 1557,
	1972052 when 1558,
	1972611 when 1559,
	1973170 when 1560,
	1973727 when 1561,
	1974283 when 1562,
	1974838 when 1563,
	1975392 when 1564,
	1975944 when 1565,
	1976496 when 1566,
	1977046 when 1567,
	1977594 when 1568,
	1978142 when 1569,
	1978688 when 1570,
	1979234 when 1571,
	1979777 when 1572,
	1980320 when 1573,
	1980862 when 1574,
	1981402 when 1575,
	1981941 when 1576,
	1982479 when 1577,
	1983015 when 1578,
	1983551 when 1579,
	1984085 when 1580,
	1984618 when 1581,
	1985149 when 1582,
	1985680 when 1583,
	1986209 when 1584,
	1986737 when 1585,
	1987264 when 1586,
	1987789 when 1587,
	1988314 when 1588,
	1988837 when 1589,
	1989359 when 1590,
	1989879 when 1591,
	1990399 when 1592,
	1990917 when 1593,
	1991434 when 1594,
	1991950 when 1595,
	1992464 when 1596,
	1992978 when 1597,
	1993490 when 1598,
	1994000 when 1599,
	1994510 when 1600,
	1995018 when 1601,
	1995526 when 1602,
	1996031 when 1603,
	1996536 when 1604,
	1997040 when 1605,
	1997542 when 1606,
	1998043 when 1607,
	1998543 when 1608,
	1999041 when 1609,
	1999538 when 1610,
	2000034 when 1611,
	2000529 when 1612,
	2001023 when 1613,
	2001515 when 1614,
	2002006 when 1615,
	2002496 when 1616,
	2002985 when 1617,
	2003472 when 1618,
	2003958 when 1619,
	2004443 when 1620,
	2004927 when 1621,
	2005409 when 1622,
	2005891 when 1623,
	2006371 when 1624,
	2006849 when 1625,
	2007327 when 1626,
	2007803 when 1627,
	2008278 when 1628,
	2008752 when 1629,
	2009224 when 1630,
	2009696 when 1631,
	2010166 when 1632,
	2010635 when 1633,
	2011102 when 1634,
	2011569 when 1635,
	2012034 when 1636,
	2012498 when 1637,
	2012960 when 1638,
	2013422 when 1639,
	2013882 when 1640,
	2014341 when 1641,
	2014798 when 1642,
	2015255 when 1643,
	2015710 when 1644,
	2016164 when 1645,
	2016617 when 1646,
	2017068 when 1647,
	2017518 when 1648,
	2017967 when 1649,
	2018415 when 1650,
	2018861 when 1651,
	2019307 when 1652,
	2019751 when 1653,
	2020193 when 1654,
	2020635 when 1655,
	2021075 when 1656,
	2021514 when 1657,
	2021952 when 1658,
	2022388 when 1659,
	2022824 when 1660,
	2023258 when 1661,
	2023690 when 1662,
	2024122 when 1663,
	2024552 when 1664,
	2024981 when 1665,
	2025409 when 1666,
	2025835 when 1667,
	2026261 when 1668,
	2026685 when 1669,
	2027107 when 1670,
	2027529 when 1671,
	2027949 when 1672,
	2028368 when 1673,
	2028786 when 1674,
	2029202 when 1675,
	2029618 when 1676,
	2030032 when 1677,
	2030444 when 1678,
	2030856 when 1679,
	2031266 when 1680,
	2031675 when 1681,
	2032083 when 1682,
	2032489 when 1683,
	2032895 when 1684,
	2033299 when 1685,
	2033701 when 1686,
	2034103 when 1687,
	2034503 when 1688,
	2034902 when 1689,
	2035300 when 1690,
	2035696 when 1691,
	2036091 when 1692,
	2036485 when 1693,
	2036878 when 1694,
	2037269 when 1695,
	2037659 when 1696,
	2038048 when 1697,
	2038436 when 1698,
	2038822 when 1699,
	2039208 when 1700,
	2039591 when 1701,
	2039974 when 1702,
	2040355 when 1703,
	2040735 when 1704,
	2041114 when 1705,
	2041492 when 1706,
	2041868 when 1707,
	2042243 when 1708,
	2042617 when 1709,
	2042990 when 1710,
	2043361 when 1711,
	2043731 when 1712,
	2044100 when 1713,
	2044467 when 1714,
	2044833 when 1715,
	2045198 when 1716,
	2045562 when 1717,
	2045925 when 1718,
	2046286 when 1719,
	2046646 when 1720,
	2047004 when 1721,
	2047362 when 1722,
	2047718 when 1723,
	2048073 when 1724,
	2048427 when 1725,
	2048779 when 1726,
	2049130 when 1727,
	2049480 when 1728,
	2049828 when 1729,
	2050176 when 1730,
	2050522 when 1731,
	2050866 when 1732,
	2051210 when 1733,
	2051552 when 1734,
	2051893 when 1735,
	2052233 when 1736,
	2052571 when 1737,
	2052909 when 1738,
	2053244 when 1739,
	2053579 when 1740,
	2053912 when 1741,
	2054245 when 1742,
	2054575 when 1743,
	2054905 when 1744,
	2055233 when 1745,
	2055560 when 1746,
	2055886 when 1747,
	2056211 when 1748,
	2056534 when 1749,
	2056856 when 1750,
	2057177 when 1751,
	2057496 when 1752,
	2057814 when 1753,
	2058131 when 1754,
	2058447 when 1755,
	2058761 when 1756,
	2059074 when 1757,
	2059386 when 1758,
	2059696 when 1759,
	2060006 when 1760,
	2060314 when 1761,
	2060620 when 1762,
	2060926 when 1763,
	2061230 when 1764,
	2061533 when 1765,
	2061835 when 1766,
	2062135 when 1767,
	2062434 when 1768,
	2062732 when 1769,
	2063028 when 1770,
	2063324 when 1771,
	2063618 when 1772,
	2063910 when 1773,
	2064202 when 1774,
	2064492 when 1775,
	2064781 when 1776,
	2065069 when 1777,
	2065355 when 1778,
	2065640 when 1779,
	2065924 when 1780,
	2066207 when 1781,
	2066488 when 1782,
	2066768 when 1783,
	2067047 when 1784,
	2067324 when 1785,
	2067600 when 1786,
	2067875 when 1787,
	2068149 when 1788,
	2068421 when 1789,
	2068692 when 1790,
	2068962 when 1791,
	2069230 when 1792,
	2069498 when 1793,
	2069764 when 1794,
	2070028 when 1795,
	2070292 when 1796,
	2070554 when 1797,
	2070815 when 1798,
	2071074 when 1799,
	2071333 when 1800,
	2071590 when 1801,
	2071845 when 1802,
	2072100 when 1803,
	2072353 when 1804,
	2072605 when 1805,
	2072856 when 1806,
	2073105 when 1807,
	2073353 when 1808,
	2073600 when 1809,
	2073845 when 1810,
	2074090 when 1811,
	2074332 when 1812,
	2074574 when 1813,
	2074815 when 1814,
	2075054 when 1815,
	2075292 when 1816,
	2075528 when 1817,
	2075763 when 1818,
	2075997 when 1819,
	2076230 when 1820,
	2076462 when 1821,
	2076692 when 1822,
	2076921 when 1823,
	2077148 when 1824,
	2077374 when 1825,
	2077600 when 1826,
	2077823 when 1827,
	2078046 when 1828,
	2078267 when 1829,
	2078487 when 1830,
	2078705 when 1831,
	2078923 when 1832,
	2079139 when 1833,
	2079354 when 1834,
	2079567 when 1835,
	2079779 when 1836,
	2079990 when 1837,
	2080200 when 1838,
	2080408 when 1839,
	2080615 when 1840,
	2080821 when 1841,
	2081026 when 1842,
	2081229 when 1843,
	2081431 when 1844,
	2081631 when 1845,
	2081831 when 1846,
	2082029 when 1847,
	2082226 when 1848,
	2082421 when 1849,
	2082616 when 1850,
	2082808 when 1851,
	2083000 when 1852,
	2083191 when 1853,
	2083380 when 1854,
	2083567 when 1855,
	2083754 when 1856,
	2083939 when 1857,
	2084123 when 1858,
	2084306 when 1859,
	2084487 when 1860,
	2084667 when 1861,
	2084846 when 1862,
	2085024 when 1863,
	2085200 when 1864,
	2085375 when 1865,
	2085549 when 1866,
	2085721 when 1867,
	2085892 when 1868,
	2086062 when 1869,
	2086230 when 1870,
	2086398 when 1871,
	2086564 when 1872,
	2086728 when 1873,
	2086892 when 1874,
	2087054 when 1875,
	2087214 when 1876,
	2087374 when 1877,
	2087532 when 1878,
	2087689 when 1879,
	2087845 when 1880,
	2087999 when 1881,
	2088152 when 1882,
	2088304 when 1883,
	2088454 when 1884,
	2088604 when 1885,
	2088752 when 1886,
	2088898 when 1887,
	2089044 when 1888,
	2089188 when 1889,
	2089330 when 1890,
	2089472 when 1891,
	2089612 when 1892,
	2089751 when 1893,
	2089889 when 1894,
	2090025 when 1895,
	2090160 when 1896,
	2090294 when 1897,
	2090426 when 1898,
	2090557 when 1899,
	2090687 when 1900,
	2090816 when 1901,
	2090943 when 1902,
	2091069 when 1903,
	2091194 when 1904,
	2091317 when 1905,
	2091439 when 1906,
	2091560 when 1907,
	2091680 when 1908,
	2091798 when 1909,
	2091915 when 1910,
	2092031 when 1911,
	2092145 when 1912,
	2092258 when 1913,
	2092370 when 1914,
	2092481 when 1915,
	2092590 when 1916,
	2092698 when 1917,
	2092804 when 1918,
	2092910 when 1919,
	2093014 when 1920,
	2093117 when 1921,
	2093218 when 1922,
	2093318 when 1923,
	2093417 when 1924,
	2093515 when 1925,
	2093611 when 1926,
	2093706 when 1927,
	2093800 when 1928,
	2093892 when 1929,
	2093983 when 1930,
	2094073 when 1931,
	2094162 when 1932,
	2094249 when 1933,
	2094335 when 1934,
	2094420 when 1935,
	2094503 when 1936,
	2094585 when 1937,
	2094666 when 1938,
	2094746 when 1939,
	2094824 when 1940,
	2094901 when 1941,
	2094976 when 1942,
	2095051 when 1943,
	2095124 when 1944,
	2095196 when 1945,
	2095266 when 1946,
	2095335 when 1947,
	2095403 when 1948,
	2095470 when 1949,
	2095535 when 1950,
	2095599 when 1951,
	2095662 when 1952,
	2095723 when 1953,
	2095783 when 1954,
	2095842 when 1955,
	2095900 when 1956,
	2095956 when 1957,
	2096011 when 1958,
	2096065 when 1959,
	2096117 when 1960,
	2096168 when 1961,
	2096218 when 1962,
	2096267 when 1963,
	2096314 when 1964,
	2096360 when 1965,
	2096404 when 1966,
	2096448 when 1967,
	2096490 when 1968,
	2096530 when 1969,
	2096570 when 1970,
	2096608 when 1971,
	2096645 when 1972,
	2096680 when 1973,
	2096715 when 1974,
	2096748 when 1975,
	2096779 when 1976,
	2096810 when 1977,
	2096839 when 1978,
	2096867 when 1979,
	2096893 when 1980,
	2096919 when 1981,
	2096942 when 1982,
	2096965 when 1983,
	2096986 when 1984,
	2097006 when 1985,
	2097025 when 1986,
	2097043 when 1987,
	2097059 when 1988,
	2097074 when 1989,
	2097087 when 1990,
	2097100 when 1991,
	2097111 when 1992,
	2097120 when 1993,
	2097129 when 1994,
	2097136 when 1995,
	2097142 when 1996,
	2097146 when 1997,
	2097149 when 1998,
	2097151 when 1999,
	2097152 when 2000,
	2097151 when 2001,
	2097149 when 2002,
	2097146 when 2003,
	2097142 when 2004,
	2097136 when 2005,
	2097129 when 2006,
	2097120 when 2007,
	2097111 when 2008,
	2097100 when 2009,
	2097087 when 2010,
	2097074 when 2011,
	2097059 when 2012,
	2097043 when 2013,
	2097025 when 2014,
	2097006 when 2015,
	2096986 when 2016,
	2096965 when 2017,
	2096942 when 2018,
	2096919 when 2019,
	2096893 when 2020,
	2096867 when 2021,
	2096839 when 2022,
	2096810 when 2023,
	2096779 when 2024,
	2096748 when 2025,
	2096715 when 2026,
	2096680 when 2027,
	2096645 when 2028,
	2096608 when 2029,
	2096570 when 2030,
	2096530 when 2031,
	2096490 when 2032,
	2096448 when 2033,
	2096404 when 2034,
	2096360 when 2035,
	2096314 when 2036,
	2096267 when 2037,
	2096218 when 2038,
	2096168 when 2039,
	2096117 when 2040,
	2096065 when 2041,
	2096011 when 2042,
	2095956 when 2043,
	2095900 when 2044,
	2095842 when 2045,
	2095783 when 2046,
	2095723 when 2047,
	2095662 when 2048,
	2095599 when 2049,
	2095535 when 2050,
	2095470 when 2051,
	2095403 when 2052,
	2095335 when 2053,
	2095266 when 2054,
	2095196 when 2055,
	2095124 when 2056,
	2095051 when 2057,
	2094976 when 2058,
	2094901 when 2059,
	2094824 when 2060,
	2094746 when 2061,
	2094666 when 2062,
	2094585 when 2063,
	2094503 when 2064,
	2094420 when 2065,
	2094335 when 2066,
	2094249 when 2067,
	2094162 when 2068,
	2094073 when 2069,
	2093983 when 2070,
	2093892 when 2071,
	2093800 when 2072,
	2093706 when 2073,
	2093611 when 2074,
	2093515 when 2075,
	2093417 when 2076,
	2093318 when 2077,
	2093218 when 2078,
	2093117 when 2079,
	2093014 when 2080,
	2092910 when 2081,
	2092804 when 2082,
	2092698 when 2083,
	2092590 when 2084,
	2092481 when 2085,
	2092370 when 2086,
	2092258 when 2087,
	2092145 when 2088,
	2092031 when 2089,
	2091915 when 2090,
	2091798 when 2091,
	2091680 when 2092,
	2091560 when 2093,
	2091439 when 2094,
	2091317 when 2095,
	2091194 when 2096,
	2091069 when 2097,
	2090943 when 2098,
	2090816 when 2099,
	2090687 when 2100,
	2090557 when 2101,
	2090426 when 2102,
	2090294 when 2103,
	2090160 when 2104,
	2090025 when 2105,
	2089889 when 2106,
	2089751 when 2107,
	2089612 when 2108,
	2089472 when 2109,
	2089330 when 2110,
	2089188 when 2111,
	2089044 when 2112,
	2088898 when 2113,
	2088752 when 2114,
	2088604 when 2115,
	2088454 when 2116,
	2088304 when 2117,
	2088152 when 2118,
	2087999 when 2119,
	2087845 when 2120,
	2087689 when 2121,
	2087532 when 2122,
	2087374 when 2123,
	2087214 when 2124,
	2087054 when 2125,
	2086892 when 2126,
	2086728 when 2127,
	2086564 when 2128,
	2086398 when 2129,
	2086230 when 2130,
	2086062 when 2131,
	2085892 when 2132,
	2085721 when 2133,
	2085549 when 2134,
	2085375 when 2135,
	2085200 when 2136,
	2085024 when 2137,
	2084846 when 2138,
	2084667 when 2139,
	2084487 when 2140,
	2084306 when 2141,
	2084123 when 2142,
	2083939 when 2143,
	2083754 when 2144,
	2083567 when 2145,
	2083380 when 2146,
	2083191 when 2147,
	2083000 when 2148,
	2082808 when 2149,
	2082616 when 2150,
	2082421 when 2151,
	2082226 when 2152,
	2082029 when 2153,
	2081831 when 2154,
	2081631 when 2155,
	2081431 when 2156,
	2081229 when 2157,
	2081026 when 2158,
	2080821 when 2159,
	2080615 when 2160,
	2080408 when 2161,
	2080200 when 2162,
	2079990 when 2163,
	2079779 when 2164,
	2079567 when 2165,
	2079354 when 2166,
	2079139 when 2167,
	2078923 when 2168,
	2078705 when 2169,
	2078487 when 2170,
	2078267 when 2171,
	2078046 when 2172,
	2077823 when 2173,
	2077600 when 2174,
	2077374 when 2175,
	2077148 when 2176,
	2076921 when 2177,
	2076692 when 2178,
	2076462 when 2179,
	2076230 when 2180,
	2075997 when 2181,
	2075763 when 2182,
	2075528 when 2183,
	2075292 when 2184,
	2075054 when 2185,
	2074815 when 2186,
	2074574 when 2187,
	2074332 when 2188,
	2074090 when 2189,
	2073845 when 2190,
	2073600 when 2191,
	2073353 when 2192,
	2073105 when 2193,
	2072856 when 2194,
	2072605 when 2195,
	2072353 when 2196,
	2072100 when 2197,
	2071845 when 2198,
	2071590 when 2199,
	2071333 when 2200,
	2071074 when 2201,
	2070815 when 2202,
	2070554 when 2203,
	2070292 when 2204,
	2070028 when 2205,
	2069764 when 2206,
	2069498 when 2207,
	2069230 when 2208,
	2068962 when 2209,
	2068692 when 2210,
	2068421 when 2211,
	2068149 when 2212,
	2067875 when 2213,
	2067600 when 2214,
	2067324 when 2215,
	2067047 when 2216,
	2066768 when 2217,
	2066488 when 2218,
	2066207 when 2219,
	2065924 when 2220,
	2065640 when 2221,
	2065355 when 2222,
	2065069 when 2223,
	2064781 when 2224,
	2064492 when 2225,
	2064202 when 2226,
	2063910 when 2227,
	2063618 when 2228,
	2063324 when 2229,
	2063028 when 2230,
	2062732 when 2231,
	2062434 when 2232,
	2062135 when 2233,
	2061835 when 2234,
	2061533 when 2235,
	2061230 when 2236,
	2060926 when 2237,
	2060620 when 2238,
	2060314 when 2239,
	2060006 when 2240,
	2059696 when 2241,
	2059386 when 2242,
	2059074 when 2243,
	2058761 when 2244,
	2058447 when 2245,
	2058131 when 2246,
	2057814 when 2247,
	2057496 when 2248,
	2057177 when 2249,
	2056856 when 2250,
	2056534 when 2251,
	2056211 when 2252,
	2055886 when 2253,
	2055560 when 2254,
	2055233 when 2255,
	2054905 when 2256,
	2054575 when 2257,
	2054245 when 2258,
	2053912 when 2259,
	2053579 when 2260,
	2053244 when 2261,
	2052909 when 2262,
	2052571 when 2263,
	2052233 when 2264,
	2051893 when 2265,
	2051552 when 2266,
	2051210 when 2267,
	2050866 when 2268,
	2050522 when 2269,
	2050176 when 2270,
	2049828 when 2271,
	2049480 when 2272,
	2049130 when 2273,
	2048779 when 2274,
	2048427 when 2275,
	2048073 when 2276,
	2047718 when 2277,
	2047362 when 2278,
	2047004 when 2279,
	2046646 when 2280,
	2046286 when 2281,
	2045925 when 2282,
	2045562 when 2283,
	2045198 when 2284,
	2044833 when 2285,
	2044467 when 2286,
	2044100 when 2287,
	2043731 when 2288,
	2043361 when 2289,
	2042990 when 2290,
	2042617 when 2291,
	2042243 when 2292,
	2041868 when 2293,
	2041492 when 2294,
	2041114 when 2295,
	2040735 when 2296,
	2040355 when 2297,
	2039974 when 2298,
	2039591 when 2299,
	2039208 when 2300,
	2038822 when 2301,
	2038436 when 2302,
	2038048 when 2303,
	2037659 when 2304,
	2037269 when 2305,
	2036878 when 2306,
	2036485 when 2307,
	2036091 when 2308,
	2035696 when 2309,
	2035300 when 2310,
	2034902 when 2311,
	2034503 when 2312,
	2034103 when 2313,
	2033701 when 2314,
	2033299 when 2315,
	2032895 when 2316,
	2032489 when 2317,
	2032083 when 2318,
	2031675 when 2319,
	2031266 when 2320,
	2030856 when 2321,
	2030444 when 2322,
	2030032 when 2323,
	2029618 when 2324,
	2029202 when 2325,
	2028786 when 2326,
	2028368 when 2327,
	2027949 when 2328,
	2027529 when 2329,
	2027107 when 2330,
	2026685 when 2331,
	2026261 when 2332,
	2025835 when 2333,
	2025409 when 2334,
	2024981 when 2335,
	2024552 when 2336,
	2024122 when 2337,
	2023690 when 2338,
	2023258 when 2339,
	2022824 when 2340,
	2022388 when 2341,
	2021952 when 2342,
	2021514 when 2343,
	2021075 when 2344,
	2020635 when 2345,
	2020193 when 2346,
	2019751 when 2347,
	2019307 when 2348,
	2018861 when 2349,
	2018415 when 2350,
	2017967 when 2351,
	2017518 when 2352,
	2017068 when 2353,
	2016617 when 2354,
	2016164 when 2355,
	2015710 when 2356,
	2015255 when 2357,
	2014798 when 2358,
	2014341 when 2359,
	2013882 when 2360,
	2013422 when 2361,
	2012960 when 2362,
	2012498 when 2363,
	2012034 when 2364,
	2011569 when 2365,
	2011102 when 2366,
	2010635 when 2367,
	2010166 when 2368,
	2009696 when 2369,
	2009224 when 2370,
	2008752 when 2371,
	2008278 when 2372,
	2007803 when 2373,
	2007327 when 2374,
	2006849 when 2375,
	2006371 when 2376,
	2005891 when 2377,
	2005409 when 2378,
	2004927 when 2379,
	2004443 when 2380,
	2003958 when 2381,
	2003472 when 2382,
	2002985 when 2383,
	2002496 when 2384,
	2002006 when 2385,
	2001515 when 2386,
	2001023 when 2387,
	2000529 when 2388,
	2000034 when 2389,
	1999538 when 2390,
	1999041 when 2391,
	1998543 when 2392,
	1998043 when 2393,
	1997542 when 2394,
	1997040 when 2395,
	1996536 when 2396,
	1996031 when 2397,
	1995526 when 2398,
	1995018 when 2399,
	1994510 when 2400,
	1994000 when 2401,
	1993490 when 2402,
	1992978 when 2403,
	1992464 when 2404,
	1991950 when 2405,
	1991434 when 2406,
	1990917 when 2407,
	1990399 when 2408,
	1989879 when 2409,
	1989359 when 2410,
	1988837 when 2411,
	1988314 when 2412,
	1987789 when 2413,
	1987264 when 2414,
	1986737 when 2415,
	1986209 when 2416,
	1985680 when 2417,
	1985149 when 2418,
	1984618 when 2419,
	1984085 when 2420,
	1983551 when 2421,
	1983015 when 2422,
	1982479 when 2423,
	1981941 when 2424,
	1981402 when 2425,
	1980862 when 2426,
	1980320 when 2427,
	1979777 when 2428,
	1979234 when 2429,
	1978688 when 2430,
	1978142 when 2431,
	1977594 when 2432,
	1977046 when 2433,
	1976496 when 2434,
	1975944 when 2435,
	1975392 when 2436,
	1974838 when 2437,
	1974283 when 2438,
	1973727 when 2439,
	1973170 when 2440,
	1972611 when 2441,
	1972052 when 2442,
	1971491 when 2443,
	1970929 when 2444,
	1970365 when 2445,
	1969800 when 2446,
	1969235 when 2447,
	1968668 when 2448,
	1968099 when 2449,
	1967530 when 2450,
	1966959 when 2451,
	1966387 when 2452,
	1965814 when 2453,
	1965240 when 2454,
	1964664 when 2455,
	1964087 when 2456,
	1963509 when 2457,
	1962930 when 2458,
	1962350 when 2459,
	1961768 when 2460,
	1961186 when 2461,
	1960601 when 2462,
	1960016 when 2463,
	1959430 when 2464,
	1958842 when 2465,
	1958253 when 2466,
	1957663 when 2467,
	1957072 when 2468,
	1956479 when 2469,
	1955886 when 2470,
	1955291 when 2471,
	1954695 when 2472,
	1954097 when 2473,
	1953499 when 2474,
	1952899 when 2475,
	1952298 when 2476,
	1951696 when 2477,
	1951093 when 2478,
	1950488 when 2479,
	1949883 when 2480,
	1949276 when 2481,
	1948668 when 2482,
	1948058 when 2483,
	1947448 when 2484,
	1946836 when 2485,
	1946223 when 2486,
	1945609 when 2487,
	1944993 when 2488,
	1944377 when 2489,
	1943759 when 2490,
	1943140 when 2491,
	1942520 when 2492,
	1941899 when 2493,
	1941276 when 2494,
	1940652 when 2495,
	1940028 when 2496,
	1939401 when 2497,
	1938774 when 2498,
	1938146 when 2499,
	1937516 when 2500,
	1936885 when 2501,
	1936253 when 2502,
	1935619 when 2503,
	1934985 when 2504,
	1934349 when 2505,
	1933712 when 2506,
	1933074 when 2507,
	1932435 when 2508,
	1931795 when 2509,
	1931153 when 2510,
	1930510 when 2511,
	1929866 when 2512,
	1929221 when 2513,
	1928574 when 2514,
	1927927 when 2515,
	1927278 when 2516,
	1926628 when 2517,
	1925977 when 2518,
	1925324 when 2519,
	1924671 when 2520,
	1924016 when 2521,
	1923360 when 2522,
	1922703 when 2523,
	1922045 when 2524,
	1921385 when 2525,
	1920725 when 2526,
	1920063 when 2527,
	1919400 when 2528,
	1918736 when 2529,
	1918070 when 2530,
	1917404 when 2531,
	1916736 when 2532,
	1916067 when 2533,
	1915397 when 2534,
	1914725 when 2535,
	1914053 when 2536,
	1913379 when 2537,
	1912704 when 2538,
	1912028 when 2539,
	1911351 when 2540,
	1910673 when 2541,
	1909993 when 2542,
	1909312 when 2543,
	1908631 when 2544,
	1907947 when 2545,
	1907263 when 2546,
	1906578 when 2547,
	1905891 when 2548,
	1905203 when 2549,
	1904514 when 2550,
	1903824 when 2551,
	1903133 when 2552,
	1902440 when 2553,
	1901747 when 2554,
	1901052 when 2555,
	1900356 when 2556,
	1899658 when 2557,
	1898960 when 2558,
	1898261 when 2559,
	1897560 when 2560,
	1896858 when 2561,
	1896155 when 2562,
	1895451 when 2563,
	1894745 when 2564,
	1894039 when 2565,
	1893331 when 2566,
	1892622 when 2567,
	1891912 when 2568,
	1891201 when 2569,
	1890488 when 2570,
	1889775 when 2571,
	1889060 when 2572,
	1888344 when 2573,
	1887627 when 2574,
	1886909 when 2575,
	1886190 when 2576,
	1885469 when 2577,
	1884747 when 2578,
	1884024 when 2579,
	1883300 when 2580,
	1882575 when 2581,
	1881849 when 2582,
	1881121 when 2583,
	1880393 when 2584,
	1879663 when 2585,
	1878932 when 2586,
	1878200 when 2587,
	1877466 when 2588,
	1876732 when 2589,
	1875996 when 2590,
	1875259 when 2591,
	1874521 when 2592,
	1873782 when 2593,
	1873042 when 2594,
	1872301 when 2595,
	1871558 when 2596,
	1870814 when 2597,
	1870069 when 2598,
	1869323 when 2599,
	1868576 when 2600,
	1867828 when 2601,
	1867078 when 2602,
	1866328 when 2603,
	1865576 when 2604,
	1864823 when 2605,
	1864069 when 2606,
	1863314 when 2607,
	1862557 when 2608,
	1861800 when 2609,
	1861041 when 2610,
	1860281 when 2611,
	1859520 when 2612,
	1858758 when 2613,
	1857995 when 2614,
	1857230 when 2615,
	1856465 when 2616,
	1855698 when 2617,
	1854930 when 2618,
	1854161 when 2619,
	1853391 when 2620,
	1852620 when 2621,
	1851847 when 2622,
	1851074 when 2623,
	1850299 when 2624,
	1849523 when 2625,
	1848746 when 2626,
	1847968 when 2627,
	1847188 when 2628,
	1846408 when 2629,
	1845627 when 2630,
	1844844 when 2631,
	1844060 when 2632,
	1843275 when 2633,
	1842489 when 2634,
	1841702 when 2635,
	1840913 when 2636,
	1840124 when 2637,
	1839333 when 2638,
	1838541 when 2639,
	1837748 when 2640,
	1836954 when 2641,
	1836159 when 2642,
	1835363 when 2643,
	1834565 when 2644,
	1833767 when 2645,
	1832967 when 2646,
	1832166 when 2647,
	1831364 when 2648,
	1830561 when 2649,
	1829757 when 2650,
	1828951 when 2651,
	1828145 when 2652,
	1827337 when 2653,
	1826528 when 2654,
	1825719 when 2655,
	1824908 when 2656,
	1824095 when 2657,
	1823282 when 2658,
	1822468 when 2659,
	1821652 when 2660,
	1820836 when 2661,
	1820018 when 2662,
	1819199 when 2663,
	1818379 when 2664,
	1817558 when 2665,
	1816736 when 2666,
	1815912 when 2667,
	1815088 when 2668,
	1814262 when 2669,
	1813436 when 2670,
	1812608 when 2671,
	1811779 when 2672,
	1810949 when 2673,
	1810117 when 2674,
	1809285 when 2675,
	1808452 when 2676,
	1807617 when 2677,
	1806782 when 2678,
	1805945 when 2679,
	1805107 when 2680,
	1804268 when 2681,
	1803428 when 2682,
	1802587 when 2683,
	1801744 when 2684,
	1800901 when 2685,
	1800056 when 2686,
	1799211 when 2687,
	1798364 when 2688,
	1797516 when 2689,
	1796667 when 2690,
	1795817 when 2691,
	1794966 when 2692,
	1794113 when 2693,
	1793260 when 2694,
	1792405 when 2695,
	1791550 when 2696,
	1790693 when 2697,
	1789835 when 2698,
	1788976 when 2699,
	1788116 when 2700,
	1787255 when 2701,
	1786393 when 2702,
	1785529 when 2703,
	1784665 when 2704,
	1783799 when 2705,
	1782933 when 2706,
	1782065 when 2707,
	1781196 when 2708,
	1780326 when 2709,
	1779455 when 2710,
	1778583 when 2711,
	1777709 when 2712,
	1776835 when 2713,
	1775960 when 2714,
	1775083 when 2715,
	1774205 when 2716,
	1773327 when 2717,
	1772447 when 2718,
	1771566 when 2719,
	1770684 when 2720,
	1769801 when 2721,
	1768917 when 2722,
	1768031 when 2723,
	1767145 when 2724,
	1766258 when 2725,
	1765369 when 2726,
	1764479 when 2727,
	1763589 when 2728,
	1762697 when 2729,
	1761804 when 2730,
	1760910 when 2731,
	1760015 when 2732,
	1759119 when 2733,
	1758221 when 2734,
	1757323 when 2735,
	1756424 when 2736,
	1755523 when 2737,
	1754622 when 2738,
	1753719 when 2739,
	1752815 when 2740,
	1751910 when 2741,
	1751004 when 2742,
	1750097 when 2743,
	1749189 when 2744,
	1748280 when 2745,
	1747370 when 2746,
	1746459 when 2747,
	1745546 when 2748,
	1744633 when 2749,
	1743718 when 2750,
	1742803 when 2751,
	1741886 when 2752,
	1740968 when 2753,
	1740049 when 2754,
	1739129 when 2755,
	1738208 when 2756,
	1737286 when 2757,
	1736363 when 2758,
	1735439 when 2759,
	1734514 when 2760,
	1733587 when 2761,
	1732660 when 2762,
	1731731 when 2763,
	1730802 when 2764,
	1729871 when 2765,
	1728940 when 2766,
	1728007 when 2767,
	1727073 when 2768,
	1726138 when 2769,
	1725202 when 2770,
	1724265 when 2771,
	1723327 when 2772,
	1722388 when 2773,
	1721448 when 2774,
	1720507 when 2775,
	1719564 when 2776,
	1718621 when 2777,
	1717676 when 2778,
	1716731 when 2779,
	1715784 when 2780,
	1714837 when 2781,
	1713888 when 2782,
	1712938 when 2783,
	1711987 when 2784,
	1711036 when 2785,
	1710083 when 2786,
	1709129 when 2787,
	1708174 when 2788,
	1707218 when 2789,
	1706261 when 2790,
	1705302 when 2791,
	1704343 when 2792,
	1703383 when 2793,
	1702422 when 2794,
	1701459 when 2795,
	1700496 when 2796,
	1699531 when 2797,
	1698566 when 2798,
	1697599 when 2799,
	1696632 when 2800,
	1695663 when 2801,
	1694693 when 2802,
	1693722 when 2803,
	1692751 when 2804,
	1691778 when 2805,
	1690804 when 2806,
	1689829 when 2807,
	1688853 when 2808,
	1687876 when 2809,
	1686898 when 2810,
	1685919 when 2811,
	1684939 when 2812,
	1683958 when 2813,
	1682975 when 2814,
	1681992 when 2815,
	1681008 when 2816,
	1680022 when 2817,
	1679036 when 2818,
	1678049 when 2819,
	1677060 when 2820,
	1676071 when 2821,
	1675080 when 2822,
	1674089 when 2823,
	1673096 when 2824,
	1672103 when 2825,
	1671108 when 2826,
	1670112 when 2827,
	1669116 when 2828,
	1668118 when 2829,
	1667119 when 2830,
	1666119 when 2831,
	1665119 when 2832,
	1664117 when 2833,
	1663114 when 2834,
	1662110 when 2835,
	1661105 when 2836,
	1660099 when 2837,
	1659092 when 2838,
	1658084 when 2839,
	1657075 when 2840,
	1656065 when 2841,
	1655054 when 2842,
	1654042 when 2843,
	1653029 when 2844,
	1652015 when 2845,
	1651000 when 2846,
	1649984 when 2847,
	1648966 when 2848,
	1647948 when 2849,
	1646929 when 2850,
	1645909 when 2851,
	1644888 when 2852,
	1643865 when 2853,
	1642842 when 2854,
	1641818 when 2855,
	1640792 when 2856,
	1639766 when 2857,
	1638739 when 2858,
	1637711 when 2859,
	1636681 when 2860,
	1635651 when 2861,
	1634619 when 2862,
	1633587 when 2863,
	1632554 when 2864,
	1631519 when 2865,
	1630484 when 2866,
	1629448 when 2867,
	1628410 when 2868,
	1627372 when 2869,
	1626332 when 2870,
	1625292 when 2871,
	1624251 when 2872,
	1623208 when 2873,
	1622165 when 2874,
	1621120 when 2875,
	1620075 when 2876,
	1619029 when 2877,
	1617981 when 2878,
	1616933 when 2879,
	1615883 when 2880,
	1614833 when 2881,
	1613782 when 2882,
	1612729 when 2883,
	1611676 when 2884,
	1610621 when 2885,
	1609566 when 2886,
	1608510 when 2887,
	1607452 when 2888,
	1606394 when 2889,
	1605335 when 2890,
	1604274 when 2891,
	1603213 when 2892,
	1602151 when 2893,
	1601087 when 2894,
	1600023 when 2895,
	1598958 when 2896,
	1597892 when 2897,
	1596824 when 2898,
	1595756 when 2899,
	1594687 when 2900,
	1593617 when 2901,
	1592546 when 2902,
	1591473 when 2903,
	1590400 when 2904,
	1589326 when 2905,
	1588251 when 2906,
	1587175 when 2907,
	1586098 when 2908,
	1585020 when 2909,
	1583941 when 2910,
	1582861 when 2911,
	1581780 when 2912,
	1580698 when 2913,
	1579615 when 2914,
	1578531 when 2915,
	1577446 when 2916,
	1576360 when 2917,
	1575273 when 2918,
	1574186 when 2919,
	1573097 when 2920,
	1572007 when 2921,
	1570916 when 2922,
	1569825 when 2923,
	1568732 when 2924,
	1567639 when 2925,
	1566544 when 2926,
	1565448 when 2927,
	1564352 when 2928,
	1563254 when 2929,
	1562156 when 2930,
	1561057 when 2931,
	1559956 when 2932,
	1558855 when 2933,
	1557753 when 2934,
	1556649 when 2935,
	1555545 when 2936,
	1554440 when 2937,
	1553334 when 2938,
	1552227 when 2939,
	1551119 when 2940,
	1550010 when 2941,
	1548900 when 2942,
	1547789 when 2943,
	1546677 when 2944,
	1545564 when 2945,
	1544451 when 2946,
	1543336 when 2947,
	1542220 when 2948,
	1541103 when 2949,
	1539986 when 2950,
	1538867 when 2951,
	1537748 when 2952,
	1536627 when 2953,
	1535506 when 2954,
	1534384 when 2955,
	1533261 when 2956,
	1532136 when 2957,
	1531011 when 2958,
	1529885 when 2959,
	1528758 when 2960,
	1527630 when 2961,
	1526501 when 2962,
	1525371 when 2963,
	1524240 when 2964,
	1523109 when 2965,
	1521976 when 2966,
	1520842 when 2967,
	1519708 when 2968,
	1518572 when 2969,
	1517436 when 2970,
	1516298 when 2971,
	1515160 when 2972,
	1514021 when 2973,
	1512881 when 2974,
	1511740 when 2975,
	1510598 when 2976,
	1509455 when 2977,
	1508311 when 2978,
	1507166 when 2979,
	1506020 when 2980,
	1504873 when 2981,
	1503726 when 2982,
	1502577 when 2983,
	1501428 when 2984,
	1500277 when 2985,
	1499126 when 2986,
	1497974 when 2987,
	1496820 when 2988,
	1495666 when 2989,
	1494511 when 2990,
	1493355 when 2991,
	1492198 when 2992,
	1491041 when 2993,
	1489882 when 2994,
	1488722 when 2995,
	1487562 when 2996,
	1486400 when 2997,
	1485238 when 2998,
	1484075 when 2999,
	1482910 when 3000,
	1481745 when 3001,
	1480579 when 3002,
	1479412 when 3003,
	1478244 when 3004,
	1477076 when 3005,
	1475906 when 3006,
	1474735 when 3007,
	1473564 when 3008,
	1472391 when 3009,
	1471218 when 3010,
	1470044 when 3011,
	1468869 when 3012,
	1467693 when 3013,
	1466516 when 3014,
	1465338 when 3015,
	1464159 when 3016,
	1462979 when 3017,
	1461799 when 3018,
	1460617 when 3019,
	1459435 when 3020,
	1458252 when 3021,
	1457067 when 3022,
	1455882 when 3023,
	1454696 when 3024,
	1453510 when 3025,
	1452322 when 3026,
	1451133 when 3027,
	1449944 when 3028,
	1448753 when 3029,
	1447562 when 3030,
	1446370 when 3031,
	1445176 when 3032,
	1443982 when 3033,
	1442787 when 3034,
	1441592 when 3035,
	1440395 when 3036,
	1439197 when 3037,
	1437999 when 3038,
	1436800 when 3039,
	1435599 when 3040,
	1434398 when 3041,
	1433196 when 3042,
	1431993 when 3043,
	1430790 when 3044,
	1429585 when 3045,
	1428379 when 3046,
	1427173 when 3047,
	1425966 when 3048,
	1424757 when 3049,
	1423548 when 3050,
	1422338 when 3051,
	1421128 when 3052,
	1419916 when 3053,
	1418703 when 3054,
	1417490 when 3055,
	1416276 when 3056,
	1415060 when 3057,
	1413844 when 3058,
	1412627 when 3059,
	1411410 when 3060,
	1410191 when 3061,
	1408971 when 3062,
	1407751 when 3063,
	1406530 when 3064,
	1405307 when 3065,
	1404084 when 3066,
	1402861 when 3067,
	1401636 when 3068,
	1400410 when 3069,
	1399184 when 3070,
	1397956 when 3071,
	1396728 when 3072,
	1395499 when 3073,
	1394269 when 3074,
	1393038 when 3075,
	1391807 when 3076,
	1390574 when 3077,
	1389341 when 3078,
	1388107 when 3079,
	1386872 when 3080,
	1385636 when 3081,
	1384399 when 3082,
	1383161 when 3083,
	1381923 when 3084,
	1380683 when 3085,
	1379443 when 3086,
	1378202 when 3087,
	1376960 when 3088,
	1375717 when 3089,
	1374474 when 3090,
	1373229 when 3091,
	1371984 when 3092,
	1370738 when 3093,
	1369491 when 3094,
	1368243 when 3095,
	1366994 when 3096,
	1365745 when 3097,
	1364495 when 3098,
	1363243 when 3099,
	1361991 when 3100,
	1360738 when 3101,
	1359485 when 3102,
	1358230 when 3103,
	1356975 when 3104,
	1355718 when 3105,
	1354461 when 3106,
	1353203 when 3107,
	1351945 when 3108,
	1350685 when 3109,
	1349425 when 3110,
	1348164 when 3111,
	1346901 when 3112,
	1345639 when 3113,
	1344375 when 3114,
	1343110 when 3115,
	1341845 when 3116,
	1340579 when 3117,
	1339312 when 3118,
	1338044 when 3119,
	1336775 when 3120,
	1335505 when 3121,
	1334235 when 3122,
	1332964 when 3123,
	1331692 when 3124,
	1330419 when 3125,
	1329146 when 3126,
	1327871 when 3127,
	1326596 when 3128,
	1325320 when 3129,
	1324043 when 3130,
	1322765 when 3131,
	1321487 when 3132,
	1320207 when 3133,
	1318927 when 3134,
	1317646 when 3135,
	1316364 when 3136,
	1315082 when 3137,
	1313798 when 3138,
	1312514 when 3139,
	1311229 when 3140,
	1309943 when 3141,
	1308656 when 3142,
	1307369 when 3143,
	1306081 when 3144,
	1304792 when 3145,
	1303502 when 3146,
	1302211 when 3147,
	1300920 when 3148,
	1299627 when 3149,
	1298334 when 3150,
	1297040 when 3151,
	1295746 when 3152,
	1294450 when 3153,
	1293154 when 3154,
	1291857 when 3155,
	1290559 when 3156,
	1289260 when 3157,
	1287961 when 3158,
	1286660 when 3159,
	1285359 when 3160,
	1284057 when 3161,
	1282755 when 3162,
	1281451 when 3163,
	1280147 when 3164,
	1278842 when 3165,
	1277536 when 3166,
	1276230 when 3167,
	1274922 when 3168,
	1273614 when 3169,
	1272305 when 3170,
	1270995 when 3171,
	1269685 when 3172,
	1268374 when 3173,
	1267061 when 3174,
	1265749 when 3175,
	1264435 when 3176,
	1263120 when 3177,
	1261805 when 3178,
	1260489 when 3179,
	1259172 when 3180,
	1257855 when 3181,
	1256537 when 3182,
	1255218 when 3183,
	1253898 when 3184,
	1252577 when 3185,
	1251256 when 3186,
	1249933 when 3187,
	1248610 when 3188,
	1247287 when 3189,
	1245962 when 3190,
	1244637 when 3191,
	1243311 when 3192,
	1241984 when 3193,
	1240656 when 3194,
	1239328 when 3195,
	1237999 when 3196,
	1236669 when 3197,
	1235339 when 3198,
	1234007 when 3199,
	1232675 when 3200,
	1231342 when 3201,
	1230008 when 3202,
	1228674 when 3203,
	1227339 when 3204,
	1226003 when 3205,
	1224666 when 3206,
	1223329 when 3207,
	1221991 when 3208,
	1220652 when 3209,
	1219312 when 3210,
	1217971 when 3211,
	1216630 when 3212,
	1215288 when 3213,
	1213945 when 3214,
	1212602 when 3215,
	1211258 when 3216,
	1209913 when 3217,
	1208567 when 3218,
	1207221 when 3219,
	1205873 when 3220,
	1204525 when 3221,
	1203177 when 3222,
	1201827 when 3223,
	1200477 when 3224,
	1199126 when 3225,
	1197775 when 3226,
	1196422 when 3227,
	1195069 when 3228,
	1193715 when 3229,
	1192361 when 3230,
	1191005 when 3231,
	1189649 when 3232,
	1188292 when 3233,
	1186935 when 3234,
	1185577 when 3235,
	1184218 when 3236,
	1182858 when 3237,
	1181497 when 3238,
	1180136 when 3239,
	1178774 when 3240,
	1177412 when 3241,
	1176048 when 3242,
	1174684 when 3243,
	1173319 when 3244,
	1171954 when 3245,
	1170588 when 3246,
	1169221 when 3247,
	1167853 when 3248,
	1166484 when 3249,
	1165115 when 3250,
	1163745 when 3251,
	1162375 when 3252,
	1161003 when 3253,
	1159631 when 3254,
	1158259 when 3255,
	1156885 when 3256,
	1155511 when 3257,
	1154136 when 3258,
	1152761 when 3259,
	1151384 when 3260,
	1150007 when 3261,
	1148630 when 3262,
	1147251 when 3263,
	1145872 when 3264,
	1144492 when 3265,
	1143112 when 3266,
	1141730 when 3267,
	1140348 when 3268,
	1138966 when 3269,
	1137582 when 3270,
	1136198 when 3271,
	1134814 when 3272,
	1133428 when 3273,
	1132042 when 3274,
	1130655 when 3275,
	1129267 when 3276,
	1127879 when 3277,
	1126490 when 3278,
	1125101 when 3279,
	1123710 when 3280,
	1122319 when 3281,
	1120927 when 3282,
	1119535 when 3283,
	1118142 when 3284,
	1116748 when 3285,
	1115354 when 3286,
	1113958 when 3287,
	1112563 when 3288,
	1111166 when 3289,
	1109769 when 3290,
	1108371 when 3291,
	1106972 when 3292,
	1105573 when 3293,
	1104173 when 3294,
	1102772 when 3295,
	1101371 when 3296,
	1099969 when 3297,
	1098566 when 3298,
	1097163 when 3299,
	1095759 when 3300,
	1094354 when 3301,
	1092949 when 3302,
	1091543 when 3303,
	1090136 when 3304,
	1088729 when 3305,
	1087320 when 3306,
	1085912 when 3307,
	1084502 when 3308,
	1083092 when 3309,
	1081681 when 3310,
	1080270 when 3311,
	1078858 when 3312,
	1077445 when 3313,
	1076032 when 3314,
	1074618 when 3315,
	1073203 when 3316,
	1071787 when 3317,
	1070371 when 3318,
	1068955 when 3319,
	1067537 when 3320,
	1066119 when 3321,
	1064700 when 3322,
	1063281 when 3323,
	1061861 when 3324,
	1060440 when 3325,
	1059019 when 3326,
	1057597 when 3327,
	1056174 when 3328,
	1054751 when 3329,
	1053327 when 3330,
	1051903 when 3331,
	1050477 when 3332,
	1049051 when 3333,
	1047625 when 3334,
	1046198 when 3335,
	1044770 when 3336,
	1043341 when 3337,
	1041912 when 3338,
	1040483 when 3339,
	1039052 when 3340,
	1037621 when 3341,
	1036189 when 3342,
	1034757 when 3343,
	1033324 when 3344,
	1031891 when 3345,
	1030456 when 3346,
	1029021 when 3347,
	1027586 when 3348,
	1026150 when 3349,
	1024713 when 3350,
	1023276 when 3351,
	1021838 when 3352,
	1020399 when 3353,
	1018960 when 3354,
	1017520 when 3355,
	1016079 when 3356,
	1014638 when 3357,
	1013196 when 3358,
	1011754 when 3359,
	1010311 when 3360,
	1008867 when 3361,
	1007423 when 3362,
	1005978 when 3363,
	1004532 when 3364,
	1003086 when 3365,
	1001639 when 3366,
	1000192 when 3367,
	998744 when 3368,
	997295 when 3369,
	995846 when 3370,
	994396 when 3371,
	992946 when 3372,
	991495 when 3373,
	990043 when 3374,
	988591 when 3375,
	987138 when 3376,
	985684 when 3377,
	984230 when 3378,
	982775 when 3379,
	981320 when 3380,
	979864 when 3381,
	978407 when 3382,
	976950 when 3383,
	975493 when 3384,
	974034 when 3385,
	972575 when 3386,
	971116 when 3387,
	969655 when 3388,
	968195 when 3389,
	966733 when 3390,
	965271 when 3391,
	963809 when 3392,
	962346 when 3393,
	960882 when 3394,
	959418 when 3395,
	957953 when 3396,
	956487 when 3397,
	955021 when 3398,
	953554 when 3399,
	952087 when 3400,
	950619 when 3401,
	949151 when 3402,
	947682 when 3403,
	946212 when 3404,
	944742 when 3405,
	943271 when 3406,
	941800 when 3407,
	940328 when 3408,
	938855 when 3409,
	937382 when 3410,
	935908 when 3411,
	934434 when 3412,
	932959 when 3413,
	931484 when 3414,
	930008 when 3415,
	928531 when 3416,
	927054 when 3417,
	925576 when 3418,
	924098 when 3419,
	922619 when 3420,
	921140 when 3421,
	919660 when 3422,
	918179 when 3423,
	916698 when 3424,
	915217 when 3425,
	913734 when 3426,
	912251 when 3427,
	910768 when 3428,
	909284 when 3429,
	907800 when 3430,
	906315 when 3431,
	904829 when 3432,
	903343 when 3433,
	901856 when 3434,
	900369 when 3435,
	898881 when 3436,
	897392 when 3437,
	895903 when 3438,
	894414 when 3439,
	892924 when 3440,
	891433 when 3441,
	889942 when 3442,
	888450 when 3443,
	886958 when 3444,
	885465 when 3445,
	883972 when 3446,
	882478 when 3447,
	880984 when 3448,
	879489 when 3449,
	877993 when 3450,
	876497 when 3451,
	875000 when 3452,
	873503 when 3453,
	872006 when 3454,
	870507 when 3455,
	869009 when 3456,
	867509 when 3457,
	866009 when 3458,
	864509 when 3459,
	863008 when 3460,
	861507 when 3461,
	860005 when 3462,
	858502 when 3463,
	856999 when 3464,
	855496 when 3465,
	853992 when 3466,
	852487 when 3467,
	850982 when 3468,
	849476 when 3469,
	847970 when 3470,
	846463 when 3471,
	844956 when 3472,
	843448 when 3473,
	841940 when 3474,
	840431 when 3475,
	838922 when 3476,
	837412 when 3477,
	835902 when 3478,
	834391 when 3479,
	832879 when 3480,
	831368 when 3481,
	829855 when 3482,
	828342 when 3483,
	826829 when 3484,
	825315 when 3485,
	823800 when 3486,
	822286 when 3487,
	820770 when 3488,
	819254 when 3489,
	817738 when 3490,
	816221 when 3491,
	814703 when 3492,
	813185 when 3493,
	811667 when 3494,
	810148 when 3495,
	808628 when 3496,
	807108 when 3497,
	805588 when 3498,
	804067 when 3499,
	802545 when 3500,
	801023 when 3501,
	799501 when 3502,
	797978 when 3503,
	796454 when 3504,
	794931 when 3505,
	793406 when 3506,
	791881 when 3507,
	790356 when 3508,
	788830 when 3509,
	787304 when 3510,
	785777 when 3511,
	784249 when 3512,
	782721 when 3513,
	781193 when 3514,
	779664 when 3515,
	778135 when 3516,
	776605 when 3517,
	775075 when 3518,
	773544 when 3519,
	772013 when 3520,
	770481 when 3521,
	768949 when 3522,
	767417 when 3523,
	765884 when 3524,
	764350 when 3525,
	762816 when 3526,
	761281 when 3527,
	759747 when 3528,
	758211 when 3529,
	756675 when 3530,
	755139 when 3531,
	753602 when 3532,
	752065 when 3533,
	750527 when 3534,
	748989 when 3535,
	747450 when 3536,
	745911 when 3537,
	744371 when 3538,
	742831 when 3539,
	741290 when 3540,
	739749 when 3541,
	738208 when 3542,
	736666 when 3543,
	735124 when 3544,
	733581 when 3545,
	732038 when 3546,
	730494 when 3547,
	728950 when 3548,
	727405 when 3549,
	725860 when 3550,
	724315 when 3551,
	722769 when 3552,
	721222 when 3553,
	719675 when 3554,
	718128 when 3555,
	716580 when 3556,
	715032 when 3557,
	713483 when 3558,
	711934 when 3559,
	710385 when 3560,
	708835 when 3561,
	707285 when 3562,
	705734 when 3563,
	704183 when 3564,
	702631 when 3565,
	701079 when 3566,
	699526 when 3567,
	697973 when 3568,
	696420 when 3569,
	694866 when 3570,
	693312 when 3571,
	691757 when 3572,
	690202 when 3573,
	688646 when 3574,
	687090 when 3575,
	685534 when 3576,
	683977 when 3577,
	682420 when 3578,
	680862 when 3579,
	679304 when 3580,
	677746 when 3581,
	676187 when 3582,
	674627 when 3583,
	673068 when 3584,
	671507 when 3585,
	669947 when 3586,
	668386 when 3587,
	666824 when 3588,
	665263 when 3589,
	663700 when 3590,
	662138 when 3591,
	660575 when 3592,
	659011 when 3593,
	657447 when 3594,
	655883 when 3595,
	654318 when 3596,
	652753 when 3597,
	651188 when 3598,
	649622 when 3599,
	648056 when 3600,
	646489 when 3601,
	644922 when 3602,
	643354 when 3603,
	641786 when 3604,
	640218 when 3605,
	638650 when 3606,
	637080 when 3607,
	635511 when 3608,
	633941 when 3609,
	632371 when 3610,
	630800 when 3611,
	629229 when 3612,
	627658 when 3613,
	626086 when 3614,
	624514 when 3615,
	622941 when 3616,
	621368 when 3617,
	619795 when 3618,
	618221 when 3619,
	616647 when 3620,
	615073 when 3621,
	613498 when 3622,
	611923 when 3623,
	610347 when 3624,
	608771 when 3625,
	607195 when 3626,
	605618 when 3627,
	604041 when 3628,
	602463 when 3629,
	600886 when 3630,
	599307 when 3631,
	597729 when 3632,
	596150 when 3633,
	594570 when 3634,
	592991 when 3635,
	591411 when 3636,
	589830 when 3637,
	588249 when 3638,
	586668 when 3639,
	585087 when 3640,
	583505 when 3641,
	581923 when 3642,
	580340 when 3643,
	578757 when 3644,
	577174 when 3645,
	575590 when 3646,
	574006 when 3647,
	572422 when 3648,
	570837 when 3649,
	569252 when 3650,
	567666 when 3651,
	566081 when 3652,
	564495 when 3653,
	562908 when 3654,
	561321 when 3655,
	559734 when 3656,
	558147 when 3657,
	556559 when 3658,
	554970 when 3659,
	553382 when 3660,
	551793 when 3661,
	550204 when 3662,
	548614 when 3663,
	547024 when 3664,
	545434 when 3665,
	543843 when 3666,
	542253 when 3667,
	540661 when 3668,
	539070 when 3669,
	537478 when 3670,
	535886 when 3671,
	534293 when 3672,
	532700 when 3673,
	531107 when 3674,
	529513 when 3675,
	527919 when 3676,
	526325 when 3677,
	524731 when 3678,
	523136 when 3679,
	521540 when 3680,
	519945 when 3681,
	518349 when 3682,
	516753 when 3683,
	515157 when 3684,
	513560 when 3685,
	511963 when 3686,
	510365 when 3687,
	508767 when 3688,
	507169 when 3689,
	505571 when 3690,
	503972 when 3691,
	502373 when 3692,
	500774 when 3693,
	499174 when 3694,
	497575 when 3695,
	495974 when 3696,
	494374 when 3697,
	492773 when 3698,
	491172 when 3699,
	489570 when 3700,
	487969 when 3701,
	486367 when 3702,
	484764 when 3703,
	483162 when 3704,
	481559 when 3705,
	479955 when 3706,
	478352 when 3707,
	476748 when 3708,
	475144 when 3709,
	473540 when 3710,
	471935 when 3711,
	470330 when 3712,
	468725 when 3713,
	467119 when 3714,
	465513 when 3715,
	463907 when 3716,
	462301 when 3717,
	460694 when 3718,
	459087 when 3719,
	457480 when 3720,
	455872 when 3721,
	454264 when 3722,
	452656 when 3723,
	451048 when 3724,
	449439 when 3725,
	447830 when 3726,
	446221 when 3727,
	444611 when 3728,
	443001 when 3729,
	441391 when 3730,
	439781 when 3731,
	438170 when 3732,
	436559 when 3733,
	434948 when 3734,
	433337 when 3735,
	431725 when 3736,
	430113 when 3737,
	428501 when 3738,
	426889 when 3739,
	425276 when 3740,
	423663 when 3741,
	422050 when 3742,
	420436 when 3743,
	418822 when 3744,
	417208 when 3745,
	415594 when 3746,
	413979 when 3747,
	412364 when 3748,
	410749 when 3749,
	409134 when 3750,
	407518 when 3751,
	405903 when 3752,
	404287 when 3753,
	402670 when 3754,
	401054 when 3755,
	399437 when 3756,
	397820 when 3757,
	396202 when 3758,
	394585 when 3759,
	392967 when 3760,
	391349 when 3761,
	389731 when 3762,
	388112 when 3763,
	386493 when 3764,
	384874 when 3765,
	383255 when 3766,
	381636 when 3767,
	380016 when 3768,
	378396 when 3769,
	376776 when 3770,
	375155 when 3771,
	373535 when 3772,
	371914 when 3773,
	370293 when 3774,
	368672 when 3775,
	367050 when 3776,
	365428 when 3777,
	363806 when 3778,
	362184 when 3779,
	360561 when 3780,
	358939 when 3781,
	357316 when 3782,
	355693 when 3783,
	354069 when 3784,
	352446 when 3785,
	350822 when 3786,
	349198 when 3787,
	347574 when 3788,
	345949 when 3789,
	344325 when 3790,
	342700 when 3791,
	341075 when 3792,
	339450 when 3793,
	337824 when 3794,
	336198 when 3795,
	334573 when 3796,
	332946 when 3797,
	331320 when 3798,
	329694 when 3799,
	328067 when 3800,
	326440 when 3801,
	324813 when 3802,
	323185 when 3803,
	321558 when 3804,
	319930 when 3805,
	318302 when 3806,
	316674 when 3807,
	315046 when 3808,
	313417 when 3809,
	311789 when 3810,
	310160 when 3811,
	308531 when 3812,
	306901 when 3813,
	305272 when 3814,
	303642 when 3815,
	302013 when 3816,
	300382 when 3817,
	298752 when 3818,
	297122 when 3819,
	295491 when 3820,
	293861 when 3821,
	292230 when 3822,
	290598 when 3823,
	288967 when 3824,
	287336 when 3825,
	285704 when 3826,
	284072 when 3827,
	282440 when 3828,
	280808 when 3829,
	279176 when 3830,
	277543 when 3831,
	275910 when 3832,
	274278 when 3833,
	272645 when 3834,
	271011 when 3835,
	269378 when 3836,
	267744 when 3837,
	266111 when 3838,
	264477 when 3839,
	262843 when 3840,
	261209 when 3841,
	259574 when 3842,
	257940 when 3843,
	256305 when 3844,
	254670 when 3845,
	253035 when 3846,
	251400 when 3847,
	249765 when 3848,
	248129 when 3849,
	246494 when 3850,
	244858 when 3851,
	243222 when 3852,
	241586 when 3853,
	239950 when 3854,
	238313 when 3855,
	236677 when 3856,
	235040 when 3857,
	233404 when 3858,
	231767 when 3859,
	230130 when 3860,
	228492 when 3861,
	226855 when 3862,
	225217 when 3863,
	223580 when 3864,
	221942 when 3865,
	220304 when 3866,
	218666 when 3867,
	217028 when 3868,
	215390 when 3869,
	213751 when 3870,
	212112 when 3871,
	210474 when 3872,
	208835 when 3873,
	207196 when 3874,
	205557 when 3875,
	203918 when 3876,
	202278 when 3877,
	200639 when 3878,
	198999 when 3879,
	197359 when 3880,
	195720 when 3881,
	194080 when 3882,
	192440 when 3883,
	190799 when 3884,
	189159 when 3885,
	187519 when 3886,
	185878 when 3887,
	184237 when 3888,
	182597 when 3889,
	180956 when 3890,
	179315 when 3891,
	177673 when 3892,
	176032 when 3893,
	174391 when 3894,
	172749 when 3895,
	171108 when 3896,
	169466 when 3897,
	167824 when 3898,
	166183 when 3899,
	164541 when 3900,
	162899 when 3901,
	161256 when 3902,
	159614 when 3903,
	157972 when 3904,
	156329 when 3905,
	154687 when 3906,
	153044 when 3907,
	151401 when 3908,
	149758 when 3909,
	148116 when 3910,
	146472 when 3911,
	144829 when 3912,
	143186 when 3913,
	141543 when 3914,
	139899 when 3915,
	138256 when 3916,
	136612 when 3917,
	134969 when 3918,
	133325 when 3919,
	131681 when 3920,
	130037 when 3921,
	128393 when 3922,
	126749 when 3923,
	125105 when 3924,
	123461 when 3925,
	121817 when 3926,
	120172 when 3927,
	118528 when 3928,
	116883 when 3929,
	115239 when 3930,
	113594 when 3931,
	111950 when 3932,
	110305 when 3933,
	108660 when 3934,
	107015 when 3935,
	105370 when 3936,
	103725 when 3937,
	102080 when 3938,
	100435 when 3939,
	98789 when 3940,
	97144 when 3941,
	95499 when 3942,
	93853 when 3943,
	92208 when 3944,
	90562 when 3945,
	88917 when 3946,
	87271 when 3947,
	85625 when 3948,
	83980 when 3949,
	82334 when 3950,
	80688 when 3951,
	79042 when 3952,
	77396 when 3953,
	75750 when 3954,
	74104 when 3955,
	72458 when 3956,
	70812 when 3957,
	69166 when 3958,
	67519 when 3959,
	65873 when 3960,
	64227 when 3961,
	62580 when 3962,
	60934 when 3963,
	59288 when 3964,
	57641 when 3965,
	55995 when 3966,
	54348 when 3967,
	52702 when 3968,
	51055 when 3969,
	49408 when 3970,
	47762 when 3971,
	46115 when 3972,
	44468 when 3973,
	42822 when 3974,
	41175 when 3975,
	39528 when 3976,
	37881 when 3977,
	36234 when 3978,
	34588 when 3979,
	32941 when 3980,
	31294 when 3981,
	29647 when 3982,
	28000 when 3983,
	26353 when 3984,
	24706 when 3985,
	23059 when 3986,
	21412 when 3987,
	19765 when 3988,
	18118 when 3989,
	16471 when 3990,
	14824 when 3991,
	13177 when 3992,
	11530 when 3993,
	9883 when 3994,
	8235 when 3995,
	6588 when 3996,
	4941 when 3997,
	3294 when 3998,
	1647 when 3999,
	0 when 4000,
	-1647 when 4001,
	-3294 when 4002,
	-4941 when 4003,
	-6588 when 4004,
	-8235 when 4005,
	-9883 when 4006,
	-11530 when 4007,
	-13177 when 4008,
	-14824 when 4009,
	-16471 when 4010,
	-18118 when 4011,
	-19765 when 4012,
	-21412 when 4013,
	-23059 when 4014,
	-24706 when 4015,
	-26353 when 4016,
	-28000 when 4017,
	-29647 when 4018,
	-31294 when 4019,
	-32941 when 4020,
	-34588 when 4021,
	-36234 when 4022,
	-37881 when 4023,
	-39528 when 4024,
	-41175 when 4025,
	-42822 when 4026,
	-44468 when 4027,
	-46115 when 4028,
	-47762 when 4029,
	-49408 when 4030,
	-51055 when 4031,
	-52702 when 4032,
	-54348 when 4033,
	-55995 when 4034,
	-57641 when 4035,
	-59288 when 4036,
	-60934 when 4037,
	-62580 when 4038,
	-64227 when 4039,
	-65873 when 4040,
	-67519 when 4041,
	-69166 when 4042,
	-70812 when 4043,
	-72458 when 4044,
	-74104 when 4045,
	-75750 when 4046,
	-77396 when 4047,
	-79042 when 4048,
	-80688 when 4049,
	-82334 when 4050,
	-83980 when 4051,
	-85625 when 4052,
	-87271 when 4053,
	-88917 when 4054,
	-90562 when 4055,
	-92208 when 4056,
	-93853 when 4057,
	-95499 when 4058,
	-97144 when 4059,
	-98789 when 4060,
	-100435 when 4061,
	-102080 when 4062,
	-103725 when 4063,
	-105370 when 4064,
	-107015 when 4065,
	-108660 when 4066,
	-110305 when 4067,
	-111950 when 4068,
	-113594 when 4069,
	-115239 when 4070,
	-116883 when 4071,
	-118528 when 4072,
	-120172 when 4073,
	-121817 when 4074,
	-123461 when 4075,
	-125105 when 4076,
	-126749 when 4077,
	-128393 when 4078,
	-130037 when 4079,
	-131681 when 4080,
	-133325 when 4081,
	-134969 when 4082,
	-136612 when 4083,
	-138256 when 4084,
	-139899 when 4085,
	-141543 when 4086,
	-143186 when 4087,
	-144829 when 4088,
	-146472 when 4089,
	-148116 when 4090,
	-149758 when 4091,
	-151401 when 4092,
	-153044 when 4093,
	-154687 when 4094,
	-156329 when 4095,
	-157972 when 4096,
	-159614 when 4097,
	-161256 when 4098,
	-162899 when 4099,
	-164541 when 4100,
	-166183 when 4101,
	-167824 when 4102,
	-169466 when 4103,
	-171108 when 4104,
	-172749 when 4105,
	-174391 when 4106,
	-176032 when 4107,
	-177673 when 4108,
	-179315 when 4109,
	-180956 when 4110,
	-182597 when 4111,
	-184237 when 4112,
	-185878 when 4113,
	-187519 when 4114,
	-189159 when 4115,
	-190799 when 4116,
	-192440 when 4117,
	-194080 when 4118,
	-195720 when 4119,
	-197359 when 4120,
	-198999 when 4121,
	-200639 when 4122,
	-202278 when 4123,
	-203918 when 4124,
	-205557 when 4125,
	-207196 when 4126,
	-208835 when 4127,
	-210474 when 4128,
	-212112 when 4129,
	-213751 when 4130,
	-215390 when 4131,
	-217028 when 4132,
	-218666 when 4133,
	-220304 when 4134,
	-221942 when 4135,
	-223580 when 4136,
	-225217 when 4137,
	-226855 when 4138,
	-228492 when 4139,
	-230130 when 4140,
	-231767 when 4141,
	-233404 when 4142,
	-235040 when 4143,
	-236677 when 4144,
	-238313 when 4145,
	-239950 when 4146,
	-241586 when 4147,
	-243222 when 4148,
	-244858 when 4149,
	-246494 when 4150,
	-248129 when 4151,
	-249765 when 4152,
	-251400 when 4153,
	-253035 when 4154,
	-254670 when 4155,
	-256305 when 4156,
	-257940 when 4157,
	-259574 when 4158,
	-261209 when 4159,
	-262843 when 4160,
	-264477 when 4161,
	-266111 when 4162,
	-267744 when 4163,
	-269378 when 4164,
	-271011 when 4165,
	-272645 when 4166,
	-274278 when 4167,
	-275910 when 4168,
	-277543 when 4169,
	-279176 when 4170,
	-280808 when 4171,
	-282440 when 4172,
	-284072 when 4173,
	-285704 when 4174,
	-287336 when 4175,
	-288967 when 4176,
	-290598 when 4177,
	-292230 when 4178,
	-293861 when 4179,
	-295491 when 4180,
	-297122 when 4181,
	-298752 when 4182,
	-300382 when 4183,
	-302013 when 4184,
	-303642 when 4185,
	-305272 when 4186,
	-306901 when 4187,
	-308531 when 4188,
	-310160 when 4189,
	-311789 when 4190,
	-313417 when 4191,
	-315046 when 4192,
	-316674 when 4193,
	-318302 when 4194,
	-319930 when 4195,
	-321558 when 4196,
	-323185 when 4197,
	-324813 when 4198,
	-326440 when 4199,
	-328067 when 4200,
	-329694 when 4201,
	-331320 when 4202,
	-332946 when 4203,
	-334573 when 4204,
	-336198 when 4205,
	-337824 when 4206,
	-339450 when 4207,
	-341075 when 4208,
	-342700 when 4209,
	-344325 when 4210,
	-345949 when 4211,
	-347574 when 4212,
	-349198 when 4213,
	-350822 when 4214,
	-352446 when 4215,
	-354069 when 4216,
	-355693 when 4217,
	-357316 when 4218,
	-358939 when 4219,
	-360561 when 4220,
	-362184 when 4221,
	-363806 when 4222,
	-365428 when 4223,
	-367050 when 4224,
	-368672 when 4225,
	-370293 when 4226,
	-371914 when 4227,
	-373535 when 4228,
	-375155 when 4229,
	-376776 when 4230,
	-378396 when 4231,
	-380016 when 4232,
	-381636 when 4233,
	-383255 when 4234,
	-384874 when 4235,
	-386493 when 4236,
	-388112 when 4237,
	-389731 when 4238,
	-391349 when 4239,
	-392967 when 4240,
	-394585 when 4241,
	-396202 when 4242,
	-397820 when 4243,
	-399437 when 4244,
	-401054 when 4245,
	-402670 when 4246,
	-404287 when 4247,
	-405903 when 4248,
	-407518 when 4249,
	-409134 when 4250,
	-410749 when 4251,
	-412364 when 4252,
	-413979 when 4253,
	-415594 when 4254,
	-417208 when 4255,
	-418822 when 4256,
	-420436 when 4257,
	-422050 when 4258,
	-423663 when 4259,
	-425276 when 4260,
	-426889 when 4261,
	-428501 when 4262,
	-430113 when 4263,
	-431725 when 4264,
	-433337 when 4265,
	-434948 when 4266,
	-436559 when 4267,
	-438170 when 4268,
	-439781 when 4269,
	-441391 when 4270,
	-443001 when 4271,
	-444611 when 4272,
	-446221 when 4273,
	-447830 when 4274,
	-449439 when 4275,
	-451048 when 4276,
	-452656 when 4277,
	-454264 when 4278,
	-455872 when 4279,
	-457480 when 4280,
	-459087 when 4281,
	-460694 when 4282,
	-462301 when 4283,
	-463907 when 4284,
	-465513 when 4285,
	-467119 when 4286,
	-468725 when 4287,
	-470330 when 4288,
	-471935 when 4289,
	-473540 when 4290,
	-475144 when 4291,
	-476748 when 4292,
	-478352 when 4293,
	-479955 when 4294,
	-481559 when 4295,
	-483162 when 4296,
	-484764 when 4297,
	-486367 when 4298,
	-487969 when 4299,
	-489570 when 4300,
	-491172 when 4301,
	-492773 when 4302,
	-494374 when 4303,
	-495974 when 4304,
	-497575 when 4305,
	-499174 when 4306,
	-500774 when 4307,
	-502373 when 4308,
	-503972 when 4309,
	-505571 when 4310,
	-507169 when 4311,
	-508767 when 4312,
	-510365 when 4313,
	-511963 when 4314,
	-513560 when 4315,
	-515157 when 4316,
	-516753 when 4317,
	-518349 when 4318,
	-519945 when 4319,
	-521540 when 4320,
	-523136 when 4321,
	-524731 when 4322,
	-526325 when 4323,
	-527919 when 4324,
	-529513 when 4325,
	-531107 when 4326,
	-532700 when 4327,
	-534293 when 4328,
	-535886 when 4329,
	-537478 when 4330,
	-539070 when 4331,
	-540661 when 4332,
	-542253 when 4333,
	-543843 when 4334,
	-545434 when 4335,
	-547024 when 4336,
	-548614 when 4337,
	-550204 when 4338,
	-551793 when 4339,
	-553382 when 4340,
	-554970 when 4341,
	-556559 when 4342,
	-558147 when 4343,
	-559734 when 4344,
	-561321 when 4345,
	-562908 when 4346,
	-564495 when 4347,
	-566081 when 4348,
	-567666 when 4349,
	-569252 when 4350,
	-570837 when 4351,
	-572422 when 4352,
	-574006 when 4353,
	-575590 when 4354,
	-577174 when 4355,
	-578757 when 4356,
	-580340 when 4357,
	-581923 when 4358,
	-583505 when 4359,
	-585087 when 4360,
	-586668 when 4361,
	-588249 when 4362,
	-589830 when 4363,
	-591411 when 4364,
	-592991 when 4365,
	-594570 when 4366,
	-596150 when 4367,
	-597729 when 4368,
	-599307 when 4369,
	-600886 when 4370,
	-602463 when 4371,
	-604041 when 4372,
	-605618 when 4373,
	-607195 when 4374,
	-608771 when 4375,
	-610347 when 4376,
	-611923 when 4377,
	-613498 when 4378,
	-615073 when 4379,
	-616647 when 4380,
	-618221 when 4381,
	-619795 when 4382,
	-621368 when 4383,
	-622941 when 4384,
	-624514 when 4385,
	-626086 when 4386,
	-627658 when 4387,
	-629229 when 4388,
	-630800 when 4389,
	-632371 when 4390,
	-633941 when 4391,
	-635511 when 4392,
	-637080 when 4393,
	-638650 when 4394,
	-640218 when 4395,
	-641786 when 4396,
	-643354 when 4397,
	-644922 when 4398,
	-646489 when 4399,
	-648056 when 4400,
	-649622 when 4401,
	-651188 when 4402,
	-652753 when 4403,
	-654318 when 4404,
	-655883 when 4405,
	-657447 when 4406,
	-659011 when 4407,
	-660575 when 4408,
	-662138 when 4409,
	-663700 when 4410,
	-665263 when 4411,
	-666824 when 4412,
	-668386 when 4413,
	-669947 when 4414,
	-671507 when 4415,
	-673068 when 4416,
	-674627 when 4417,
	-676187 when 4418,
	-677746 when 4419,
	-679304 when 4420,
	-680862 when 4421,
	-682420 when 4422,
	-683977 when 4423,
	-685534 when 4424,
	-687090 when 4425,
	-688646 when 4426,
	-690202 when 4427,
	-691757 when 4428,
	-693312 when 4429,
	-694866 when 4430,
	-696420 when 4431,
	-697973 when 4432,
	-699526 when 4433,
	-701079 when 4434,
	-702631 when 4435,
	-704183 when 4436,
	-705734 when 4437,
	-707285 when 4438,
	-708835 when 4439,
	-710385 when 4440,
	-711934 when 4441,
	-713483 when 4442,
	-715032 when 4443,
	-716580 when 4444,
	-718128 when 4445,
	-719675 when 4446,
	-721222 when 4447,
	-722769 when 4448,
	-724315 when 4449,
	-725860 when 4450,
	-727405 when 4451,
	-728950 when 4452,
	-730494 when 4453,
	-732038 when 4454,
	-733581 when 4455,
	-735124 when 4456,
	-736666 when 4457,
	-738208 when 4458,
	-739749 when 4459,
	-741290 when 4460,
	-742831 when 4461,
	-744371 when 4462,
	-745911 when 4463,
	-747450 when 4464,
	-748989 when 4465,
	-750527 when 4466,
	-752065 when 4467,
	-753602 when 4468,
	-755139 when 4469,
	-756675 when 4470,
	-758211 when 4471,
	-759747 when 4472,
	-761281 when 4473,
	-762816 when 4474,
	-764350 when 4475,
	-765884 when 4476,
	-767417 when 4477,
	-768949 when 4478,
	-770481 when 4479,
	-772013 when 4480,
	-773544 when 4481,
	-775075 when 4482,
	-776605 when 4483,
	-778135 when 4484,
	-779664 when 4485,
	-781193 when 4486,
	-782721 when 4487,
	-784249 when 4488,
	-785777 when 4489,
	-787304 when 4490,
	-788830 when 4491,
	-790356 when 4492,
	-791881 when 4493,
	-793406 when 4494,
	-794931 when 4495,
	-796454 when 4496,
	-797978 when 4497,
	-799501 when 4498,
	-801023 when 4499,
	-802545 when 4500,
	-804067 when 4501,
	-805588 when 4502,
	-807108 when 4503,
	-808628 when 4504,
	-810148 when 4505,
	-811667 when 4506,
	-813185 when 4507,
	-814703 when 4508,
	-816221 when 4509,
	-817738 when 4510,
	-819254 when 4511,
	-820770 when 4512,
	-822286 when 4513,
	-823800 when 4514,
	-825315 when 4515,
	-826829 when 4516,
	-828342 when 4517,
	-829855 when 4518,
	-831368 when 4519,
	-832879 when 4520,
	-834391 when 4521,
	-835902 when 4522,
	-837412 when 4523,
	-838922 when 4524,
	-840431 when 4525,
	-841940 when 4526,
	-843448 when 4527,
	-844956 when 4528,
	-846463 when 4529,
	-847970 when 4530,
	-849476 when 4531,
	-850982 when 4532,
	-852487 when 4533,
	-853992 when 4534,
	-855496 when 4535,
	-856999 when 4536,
	-858502 when 4537,
	-860005 when 4538,
	-861507 when 4539,
	-863008 when 4540,
	-864509 when 4541,
	-866009 when 4542,
	-867509 when 4543,
	-869009 when 4544,
	-870507 when 4545,
	-872006 when 4546,
	-873503 when 4547,
	-875000 when 4548,
	-876497 when 4549,
	-877993 when 4550,
	-879489 when 4551,
	-880984 when 4552,
	-882478 when 4553,
	-883972 when 4554,
	-885465 when 4555,
	-886958 when 4556,
	-888450 when 4557,
	-889942 when 4558,
	-891433 when 4559,
	-892924 when 4560,
	-894414 when 4561,
	-895903 when 4562,
	-897392 when 4563,
	-898881 when 4564,
	-900369 when 4565,
	-901856 when 4566,
	-903343 when 4567,
	-904829 when 4568,
	-906315 when 4569,
	-907800 when 4570,
	-909284 when 4571,
	-910768 when 4572,
	-912251 when 4573,
	-913734 when 4574,
	-915217 when 4575,
	-916698 when 4576,
	-918179 when 4577,
	-919660 when 4578,
	-921140 when 4579,
	-922619 when 4580,
	-924098 when 4581,
	-925576 when 4582,
	-927054 when 4583,
	-928531 when 4584,
	-930008 when 4585,
	-931484 when 4586,
	-932959 when 4587,
	-934434 when 4588,
	-935908 when 4589,
	-937382 when 4590,
	-938855 when 4591,
	-940328 when 4592,
	-941800 when 4593,
	-943271 when 4594,
	-944742 when 4595,
	-946212 when 4596,
	-947682 when 4597,
	-949151 when 4598,
	-950619 when 4599,
	-952087 when 4600,
	-953554 when 4601,
	-955021 when 4602,
	-956487 when 4603,
	-957953 when 4604,
	-959418 when 4605,
	-960882 when 4606,
	-962346 when 4607,
	-963809 when 4608,
	-965271 when 4609,
	-966733 when 4610,
	-968195 when 4611,
	-969655 when 4612,
	-971116 when 4613,
	-972575 when 4614,
	-974034 when 4615,
	-975493 when 4616,
	-976950 when 4617,
	-978407 when 4618,
	-979864 when 4619,
	-981320 when 4620,
	-982775 when 4621,
	-984230 when 4622,
	-985684 when 4623,
	-987138 when 4624,
	-988591 when 4625,
	-990043 when 4626,
	-991495 when 4627,
	-992946 when 4628,
	-994396 when 4629,
	-995846 when 4630,
	-997295 when 4631,
	-998744 when 4632,
	-1000192 when 4633,
	-1001639 when 4634,
	-1003086 when 4635,
	-1004532 when 4636,
	-1005978 when 4637,
	-1007423 when 4638,
	-1008867 when 4639,
	-1010311 when 4640,
	-1011754 when 4641,
	-1013196 when 4642,
	-1014638 when 4643,
	-1016079 when 4644,
	-1017520 when 4645,
	-1018960 when 4646,
	-1020399 when 4647,
	-1021838 when 4648,
	-1023276 when 4649,
	-1024713 when 4650,
	-1026150 when 4651,
	-1027586 when 4652,
	-1029021 when 4653,
	-1030456 when 4654,
	-1031891 when 4655,
	-1033324 when 4656,
	-1034757 when 4657,
	-1036189 when 4658,
	-1037621 when 4659,
	-1039052 when 4660,
	-1040483 when 4661,
	-1041912 when 4662,
	-1043341 when 4663,
	-1044770 when 4664,
	-1046198 when 4665,
	-1047625 when 4666,
	-1049051 when 4667,
	-1050477 when 4668,
	-1051903 when 4669,
	-1053327 when 4670,
	-1054751 when 4671,
	-1056174 when 4672,
	-1057597 when 4673,
	-1059019 when 4674,
	-1060440 when 4675,
	-1061861 when 4676,
	-1063281 when 4677,
	-1064700 when 4678,
	-1066119 when 4679,
	-1067537 when 4680,
	-1068955 when 4681,
	-1070371 when 4682,
	-1071787 when 4683,
	-1073203 when 4684,
	-1074618 when 4685,
	-1076032 when 4686,
	-1077445 when 4687,
	-1078858 when 4688,
	-1080270 when 4689,
	-1081681 when 4690,
	-1083092 when 4691,
	-1084502 when 4692,
	-1085912 when 4693,
	-1087320 when 4694,
	-1088729 when 4695,
	-1090136 when 4696,
	-1091543 when 4697,
	-1092949 when 4698,
	-1094354 when 4699,
	-1095759 when 4700,
	-1097163 when 4701,
	-1098566 when 4702,
	-1099969 when 4703,
	-1101371 when 4704,
	-1102772 when 4705,
	-1104173 when 4706,
	-1105573 when 4707,
	-1106972 when 4708,
	-1108371 when 4709,
	-1109769 when 4710,
	-1111166 when 4711,
	-1112563 when 4712,
	-1113958 when 4713,
	-1115354 when 4714,
	-1116748 when 4715,
	-1118142 when 4716,
	-1119535 when 4717,
	-1120927 when 4718,
	-1122319 when 4719,
	-1123710 when 4720,
	-1125101 when 4721,
	-1126490 when 4722,
	-1127879 when 4723,
	-1129267 when 4724,
	-1130655 when 4725,
	-1132042 when 4726,
	-1133428 when 4727,
	-1134814 when 4728,
	-1136198 when 4729,
	-1137582 when 4730,
	-1138966 when 4731,
	-1140348 when 4732,
	-1141730 when 4733,
	-1143112 when 4734,
	-1144492 when 4735,
	-1145872 when 4736,
	-1147251 when 4737,
	-1148630 when 4738,
	-1150007 when 4739,
	-1151384 when 4740,
	-1152761 when 4741,
	-1154136 when 4742,
	-1155511 when 4743,
	-1156885 when 4744,
	-1158259 when 4745,
	-1159631 when 4746,
	-1161003 when 4747,
	-1162375 when 4748,
	-1163745 when 4749,
	-1165115 when 4750,
	-1166484 when 4751,
	-1167853 when 4752,
	-1169221 when 4753,
	-1170588 when 4754,
	-1171954 when 4755,
	-1173319 when 4756,
	-1174684 when 4757,
	-1176048 when 4758,
	-1177412 when 4759,
	-1178774 when 4760,
	-1180136 when 4761,
	-1181497 when 4762,
	-1182858 when 4763,
	-1184218 when 4764,
	-1185577 when 4765,
	-1186935 when 4766,
	-1188292 when 4767,
	-1189649 when 4768,
	-1191005 when 4769,
	-1192361 when 4770,
	-1193715 when 4771,
	-1195069 when 4772,
	-1196422 when 4773,
	-1197775 when 4774,
	-1199126 when 4775,
	-1200477 when 4776,
	-1201827 when 4777,
	-1203177 when 4778,
	-1204525 when 4779,
	-1205873 when 4780,
	-1207221 when 4781,
	-1208567 when 4782,
	-1209913 when 4783,
	-1211258 when 4784,
	-1212602 when 4785,
	-1213945 when 4786,
	-1215288 when 4787,
	-1216630 when 4788,
	-1217971 when 4789,
	-1219312 when 4790,
	-1220652 when 4791,
	-1221991 when 4792,
	-1223329 when 4793,
	-1224666 when 4794,
	-1226003 when 4795,
	-1227339 when 4796,
	-1228674 when 4797,
	-1230008 when 4798,
	-1231342 when 4799,
	-1232675 when 4800,
	-1234007 when 4801,
	-1235339 when 4802,
	-1236669 when 4803,
	-1237999 when 4804,
	-1239328 when 4805,
	-1240656 when 4806,
	-1241984 when 4807,
	-1243311 when 4808,
	-1244637 when 4809,
	-1245962 when 4810,
	-1247287 when 4811,
	-1248610 when 4812,
	-1249933 when 4813,
	-1251256 when 4814,
	-1252577 when 4815,
	-1253898 when 4816,
	-1255218 when 4817,
	-1256537 when 4818,
	-1257855 when 4819,
	-1259172 when 4820,
	-1260489 when 4821,
	-1261805 when 4822,
	-1263120 when 4823,
	-1264435 when 4824,
	-1265749 when 4825,
	-1267061 when 4826,
	-1268374 when 4827,
	-1269685 when 4828,
	-1270995 when 4829,
	-1272305 when 4830,
	-1273614 when 4831,
	-1274922 when 4832,
	-1276230 when 4833,
	-1277536 when 4834,
	-1278842 when 4835,
	-1280147 when 4836,
	-1281451 when 4837,
	-1282755 when 4838,
	-1284057 when 4839,
	-1285359 when 4840,
	-1286660 when 4841,
	-1287961 when 4842,
	-1289260 when 4843,
	-1290559 when 4844,
	-1291857 when 4845,
	-1293154 when 4846,
	-1294450 when 4847,
	-1295746 when 4848,
	-1297040 when 4849,
	-1298334 when 4850,
	-1299627 when 4851,
	-1300920 when 4852,
	-1302211 when 4853,
	-1303502 when 4854,
	-1304792 when 4855,
	-1306081 when 4856,
	-1307369 when 4857,
	-1308656 when 4858,
	-1309943 when 4859,
	-1311229 when 4860,
	-1312514 when 4861,
	-1313798 when 4862,
	-1315082 when 4863,
	-1316364 when 4864,
	-1317646 when 4865,
	-1318927 when 4866,
	-1320207 when 4867,
	-1321487 when 4868,
	-1322765 when 4869,
	-1324043 when 4870,
	-1325320 when 4871,
	-1326596 when 4872,
	-1327871 when 4873,
	-1329146 when 4874,
	-1330419 when 4875,
	-1331692 when 4876,
	-1332964 when 4877,
	-1334235 when 4878,
	-1335505 when 4879,
	-1336775 when 4880,
	-1338044 when 4881,
	-1339312 when 4882,
	-1340579 when 4883,
	-1341845 when 4884,
	-1343110 when 4885,
	-1344375 when 4886,
	-1345639 when 4887,
	-1346901 when 4888,
	-1348164 when 4889,
	-1349425 when 4890,
	-1350685 when 4891,
	-1351945 when 4892,
	-1353203 when 4893,
	-1354461 when 4894,
	-1355718 when 4895,
	-1356975 when 4896,
	-1358230 when 4897,
	-1359485 when 4898,
	-1360738 when 4899,
	-1361991 when 4900,
	-1363243 when 4901,
	-1364495 when 4902,
	-1365745 when 4903,
	-1366994 when 4904,
	-1368243 when 4905,
	-1369491 when 4906,
	-1370738 when 4907,
	-1371984 when 4908,
	-1373229 when 4909,
	-1374474 when 4910,
	-1375717 when 4911,
	-1376960 when 4912,
	-1378202 when 4913,
	-1379443 when 4914,
	-1380683 when 4915,
	-1381923 when 4916,
	-1383161 when 4917,
	-1384399 when 4918,
	-1385636 when 4919,
	-1386872 when 4920,
	-1388107 when 4921,
	-1389341 when 4922,
	-1390574 when 4923,
	-1391807 when 4924,
	-1393038 when 4925,
	-1394269 when 4926,
	-1395499 when 4927,
	-1396728 when 4928,
	-1397956 when 4929,
	-1399184 when 4930,
	-1400410 when 4931,
	-1401636 when 4932,
	-1402861 when 4933,
	-1404084 when 4934,
	-1405307 when 4935,
	-1406530 when 4936,
	-1407751 when 4937,
	-1408971 when 4938,
	-1410191 when 4939,
	-1411410 when 4940,
	-1412627 when 4941,
	-1413844 when 4942,
	-1415060 when 4943,
	-1416276 when 4944,
	-1417490 when 4945,
	-1418703 when 4946,
	-1419916 when 4947,
	-1421128 when 4948,
	-1422338 when 4949,
	-1423548 when 4950,
	-1424757 when 4951,
	-1425966 when 4952,
	-1427173 when 4953,
	-1428379 when 4954,
	-1429585 when 4955,
	-1430790 when 4956,
	-1431993 when 4957,
	-1433196 when 4958,
	-1434398 when 4959,
	-1435599 when 4960,
	-1436800 when 4961,
	-1437999 when 4962,
	-1439197 when 4963,
	-1440395 when 4964,
	-1441592 when 4965,
	-1442787 when 4966,
	-1443982 when 4967,
	-1445176 when 4968,
	-1446370 when 4969,
	-1447562 when 4970,
	-1448753 when 4971,
	-1449944 when 4972,
	-1451133 when 4973,
	-1452322 when 4974,
	-1453510 when 4975,
	-1454696 when 4976,
	-1455882 when 4977,
	-1457067 when 4978,
	-1458252 when 4979,
	-1459435 when 4980,
	-1460617 when 4981,
	-1461799 when 4982,
	-1462979 when 4983,
	-1464159 when 4984,
	-1465338 when 4985,
	-1466516 when 4986,
	-1467693 when 4987,
	-1468869 when 4988,
	-1470044 when 4989,
	-1471218 when 4990,
	-1472391 when 4991,
	-1473564 when 4992,
	-1474735 when 4993,
	-1475906 when 4994,
	-1477076 when 4995,
	-1478244 when 4996,
	-1479412 when 4997,
	-1480579 when 4998,
	-1481745 when 4999,
	-1482910 when 5000,
	-1484075 when 5001,
	-1485238 when 5002,
	-1486400 when 5003,
	-1487562 when 5004,
	-1488722 when 5005,
	-1489882 when 5006,
	-1491041 when 5007,
	-1492198 when 5008,
	-1493355 when 5009,
	-1494511 when 5010,
	-1495666 when 5011,
	-1496820 when 5012,
	-1497974 when 5013,
	-1499126 when 5014,
	-1500277 when 5015,
	-1501428 when 5016,
	-1502577 when 5017,
	-1503726 when 5018,
	-1504873 when 5019,
	-1506020 when 5020,
	-1507166 when 5021,
	-1508311 when 5022,
	-1509455 when 5023,
	-1510598 when 5024,
	-1511740 when 5025,
	-1512881 when 5026,
	-1514021 when 5027,
	-1515160 when 5028,
	-1516298 when 5029,
	-1517436 when 5030,
	-1518572 when 5031,
	-1519708 when 5032,
	-1520842 when 5033,
	-1521976 when 5034,
	-1523109 when 5035,
	-1524240 when 5036,
	-1525371 when 5037,
	-1526501 when 5038,
	-1527630 when 5039,
	-1528758 when 5040,
	-1529885 when 5041,
	-1531011 when 5042,
	-1532136 when 5043,
	-1533261 when 5044,
	-1534384 when 5045,
	-1535506 when 5046,
	-1536627 when 5047,
	-1537748 when 5048,
	-1538867 when 5049,
	-1539986 when 5050,
	-1541103 when 5051,
	-1542220 when 5052,
	-1543336 when 5053,
	-1544451 when 5054,
	-1545564 when 5055,
	-1546677 when 5056,
	-1547789 when 5057,
	-1548900 when 5058,
	-1550010 when 5059,
	-1551119 when 5060,
	-1552227 when 5061,
	-1553334 when 5062,
	-1554440 when 5063,
	-1555545 when 5064,
	-1556649 when 5065,
	-1557753 when 5066,
	-1558855 when 5067,
	-1559956 when 5068,
	-1561057 when 5069,
	-1562156 when 5070,
	-1563254 when 5071,
	-1564352 when 5072,
	-1565448 when 5073,
	-1566544 when 5074,
	-1567639 when 5075,
	-1568732 when 5076,
	-1569825 when 5077,
	-1570916 when 5078,
	-1572007 when 5079,
	-1573097 when 5080,
	-1574186 when 5081,
	-1575273 when 5082,
	-1576360 when 5083,
	-1577446 when 5084,
	-1578531 when 5085,
	-1579615 when 5086,
	-1580698 when 5087,
	-1581780 when 5088,
	-1582861 when 5089,
	-1583941 when 5090,
	-1585020 when 5091,
	-1586098 when 5092,
	-1587175 when 5093,
	-1588251 when 5094,
	-1589326 when 5095,
	-1590400 when 5096,
	-1591473 when 5097,
	-1592546 when 5098,
	-1593617 when 5099,
	-1594687 when 5100,
	-1595756 when 5101,
	-1596824 when 5102,
	-1597892 when 5103,
	-1598958 when 5104,
	-1600023 when 5105,
	-1601087 when 5106,
	-1602151 when 5107,
	-1603213 when 5108,
	-1604274 when 5109,
	-1605335 when 5110,
	-1606394 when 5111,
	-1607452 when 5112,
	-1608510 when 5113,
	-1609566 when 5114,
	-1610621 when 5115,
	-1611676 when 5116,
	-1612729 when 5117,
	-1613782 when 5118,
	-1614833 when 5119,
	-1615883 when 5120,
	-1616933 when 5121,
	-1617981 when 5122,
	-1619029 when 5123,
	-1620075 when 5124,
	-1621120 when 5125,
	-1622165 when 5126,
	-1623208 when 5127,
	-1624251 when 5128,
	-1625292 when 5129,
	-1626332 when 5130,
	-1627372 when 5131,
	-1628410 when 5132,
	-1629448 when 5133,
	-1630484 when 5134,
	-1631519 when 5135,
	-1632554 when 5136,
	-1633587 when 5137,
	-1634619 when 5138,
	-1635651 when 5139,
	-1636681 when 5140,
	-1637711 when 5141,
	-1638739 when 5142,
	-1639766 when 5143,
	-1640792 when 5144,
	-1641818 when 5145,
	-1642842 when 5146,
	-1643865 when 5147,
	-1644888 when 5148,
	-1645909 when 5149,
	-1646929 when 5150,
	-1647948 when 5151,
	-1648966 when 5152,
	-1649984 when 5153,
	-1651000 when 5154,
	-1652015 when 5155,
	-1653029 when 5156,
	-1654042 when 5157,
	-1655054 when 5158,
	-1656065 when 5159,
	-1657075 when 5160,
	-1658084 when 5161,
	-1659092 when 5162,
	-1660099 when 5163,
	-1661105 when 5164,
	-1662110 when 5165,
	-1663114 when 5166,
	-1664117 when 5167,
	-1665119 when 5168,
	-1666119 when 5169,
	-1667119 when 5170,
	-1668118 when 5171,
	-1669116 when 5172,
	-1670112 when 5173,
	-1671108 when 5174,
	-1672103 when 5175,
	-1673096 when 5176,
	-1674089 when 5177,
	-1675080 when 5178,
	-1676071 when 5179,
	-1677060 when 5180,
	-1678049 when 5181,
	-1679036 when 5182,
	-1680022 when 5183,
	-1681008 when 5184,
	-1681992 when 5185,
	-1682975 when 5186,
	-1683958 when 5187,
	-1684939 when 5188,
	-1685919 when 5189,
	-1686898 when 5190,
	-1687876 when 5191,
	-1688853 when 5192,
	-1689829 when 5193,
	-1690804 when 5194,
	-1691778 when 5195,
	-1692751 when 5196,
	-1693722 when 5197,
	-1694693 when 5198,
	-1695663 when 5199,
	-1696632 when 5200,
	-1697599 when 5201,
	-1698566 when 5202,
	-1699531 when 5203,
	-1700496 when 5204,
	-1701459 when 5205,
	-1702422 when 5206,
	-1703383 when 5207,
	-1704343 when 5208,
	-1705302 when 5209,
	-1706261 when 5210,
	-1707218 when 5211,
	-1708174 when 5212,
	-1709129 when 5213,
	-1710083 when 5214,
	-1711036 when 5215,
	-1711987 when 5216,
	-1712938 when 5217,
	-1713888 when 5218,
	-1714837 when 5219,
	-1715784 when 5220,
	-1716731 when 5221,
	-1717676 when 5222,
	-1718621 when 5223,
	-1719564 when 5224,
	-1720507 when 5225,
	-1721448 when 5226,
	-1722388 when 5227,
	-1723327 when 5228,
	-1724265 when 5229,
	-1725202 when 5230,
	-1726138 when 5231,
	-1727073 when 5232,
	-1728007 when 5233,
	-1728940 when 5234,
	-1729871 when 5235,
	-1730802 when 5236,
	-1731731 when 5237,
	-1732660 when 5238,
	-1733587 when 5239,
	-1734514 when 5240,
	-1735439 when 5241,
	-1736363 when 5242,
	-1737286 when 5243,
	-1738208 when 5244,
	-1739129 when 5245,
	-1740049 when 5246,
	-1740968 when 5247,
	-1741886 when 5248,
	-1742803 when 5249,
	-1743718 when 5250,
	-1744633 when 5251,
	-1745546 when 5252,
	-1746459 when 5253,
	-1747370 when 5254,
	-1748280 when 5255,
	-1749189 when 5256,
	-1750097 when 5257,
	-1751004 when 5258,
	-1751910 when 5259,
	-1752815 when 5260,
	-1753719 when 5261,
	-1754622 when 5262,
	-1755523 when 5263,
	-1756424 when 5264,
	-1757323 when 5265,
	-1758221 when 5266,
	-1759119 when 5267,
	-1760015 when 5268,
	-1760910 when 5269,
	-1761804 when 5270,
	-1762697 when 5271,
	-1763589 when 5272,
	-1764479 when 5273,
	-1765369 when 5274,
	-1766258 when 5275,
	-1767145 when 5276,
	-1768031 when 5277,
	-1768917 when 5278,
	-1769801 when 5279,
	-1770684 when 5280,
	-1771566 when 5281,
	-1772447 when 5282,
	-1773327 when 5283,
	-1774205 when 5284,
	-1775083 when 5285,
	-1775960 when 5286,
	-1776835 when 5287,
	-1777709 when 5288,
	-1778583 when 5289,
	-1779455 when 5290,
	-1780326 when 5291,
	-1781196 when 5292,
	-1782065 when 5293,
	-1782933 when 5294,
	-1783799 when 5295,
	-1784665 when 5296,
	-1785529 when 5297,
	-1786393 when 5298,
	-1787255 when 5299,
	-1788116 when 5300,
	-1788976 when 5301,
	-1789835 when 5302,
	-1790693 when 5303,
	-1791550 when 5304,
	-1792405 when 5305,
	-1793260 when 5306,
	-1794113 when 5307,
	-1794966 when 5308,
	-1795817 when 5309,
	-1796667 when 5310,
	-1797516 when 5311,
	-1798364 when 5312,
	-1799211 when 5313,
	-1800056 when 5314,
	-1800901 when 5315,
	-1801744 when 5316,
	-1802587 when 5317,
	-1803428 when 5318,
	-1804268 when 5319,
	-1805107 when 5320,
	-1805945 when 5321,
	-1806782 when 5322,
	-1807617 when 5323,
	-1808452 when 5324,
	-1809285 when 5325,
	-1810117 when 5326,
	-1810949 when 5327,
	-1811779 when 5328,
	-1812608 when 5329,
	-1813436 when 5330,
	-1814262 when 5331,
	-1815088 when 5332,
	-1815912 when 5333,
	-1816736 when 5334,
	-1817558 when 5335,
	-1818379 when 5336,
	-1819199 when 5337,
	-1820018 when 5338,
	-1820836 when 5339,
	-1821652 when 5340,
	-1822468 when 5341,
	-1823282 when 5342,
	-1824095 when 5343,
	-1824908 when 5344,
	-1825719 when 5345,
	-1826528 when 5346,
	-1827337 when 5347,
	-1828145 when 5348,
	-1828951 when 5349,
	-1829757 when 5350,
	-1830561 when 5351,
	-1831364 when 5352,
	-1832166 when 5353,
	-1832967 when 5354,
	-1833767 when 5355,
	-1834565 when 5356,
	-1835363 when 5357,
	-1836159 when 5358,
	-1836954 when 5359,
	-1837748 when 5360,
	-1838541 when 5361,
	-1839333 when 5362,
	-1840124 when 5363,
	-1840913 when 5364,
	-1841702 when 5365,
	-1842489 when 5366,
	-1843275 when 5367,
	-1844060 when 5368,
	-1844844 when 5369,
	-1845627 when 5370,
	-1846408 when 5371,
	-1847188 when 5372,
	-1847968 when 5373,
	-1848746 when 5374,
	-1849523 when 5375,
	-1850299 when 5376,
	-1851074 when 5377,
	-1851847 when 5378,
	-1852620 when 5379,
	-1853391 when 5380,
	-1854161 when 5381,
	-1854930 when 5382,
	-1855698 when 5383,
	-1856465 when 5384,
	-1857230 when 5385,
	-1857995 when 5386,
	-1858758 when 5387,
	-1859520 when 5388,
	-1860281 when 5389,
	-1861041 when 5390,
	-1861800 when 5391,
	-1862557 when 5392,
	-1863314 when 5393,
	-1864069 when 5394,
	-1864823 when 5395,
	-1865576 when 5396,
	-1866328 when 5397,
	-1867078 when 5398,
	-1867828 when 5399,
	-1868576 when 5400,
	-1869323 when 5401,
	-1870069 when 5402,
	-1870814 when 5403,
	-1871558 when 5404,
	-1872301 when 5405,
	-1873042 when 5406,
	-1873782 when 5407,
	-1874521 when 5408,
	-1875259 when 5409,
	-1875996 when 5410,
	-1876732 when 5411,
	-1877466 when 5412,
	-1878200 when 5413,
	-1878932 when 5414,
	-1879663 when 5415,
	-1880393 when 5416,
	-1881121 when 5417,
	-1881849 when 5418,
	-1882575 when 5419,
	-1883300 when 5420,
	-1884024 when 5421,
	-1884747 when 5422,
	-1885469 when 5423,
	-1886190 when 5424,
	-1886909 when 5425,
	-1887627 when 5426,
	-1888344 when 5427,
	-1889060 when 5428,
	-1889775 when 5429,
	-1890488 when 5430,
	-1891201 when 5431,
	-1891912 when 5432,
	-1892622 when 5433,
	-1893331 when 5434,
	-1894039 when 5435,
	-1894745 when 5436,
	-1895451 when 5437,
	-1896155 when 5438,
	-1896858 when 5439,
	-1897560 when 5440,
	-1898261 when 5441,
	-1898960 when 5442,
	-1899658 when 5443,
	-1900356 when 5444,
	-1901052 when 5445,
	-1901747 when 5446,
	-1902440 when 5447,
	-1903133 when 5448,
	-1903824 when 5449,
	-1904514 when 5450,
	-1905203 when 5451,
	-1905891 when 5452,
	-1906578 when 5453,
	-1907263 when 5454,
	-1907947 when 5455,
	-1908631 when 5456,
	-1909312 when 5457,
	-1909993 when 5458,
	-1910673 when 5459,
	-1911351 when 5460,
	-1912028 when 5461,
	-1912704 when 5462,
	-1913379 when 5463,
	-1914053 when 5464,
	-1914725 when 5465,
	-1915397 when 5466,
	-1916067 when 5467,
	-1916736 when 5468,
	-1917404 when 5469,
	-1918070 when 5470,
	-1918736 when 5471,
	-1919400 when 5472,
	-1920063 when 5473,
	-1920725 when 5474,
	-1921385 when 5475,
	-1922045 when 5476,
	-1922703 when 5477,
	-1923360 when 5478,
	-1924016 when 5479,
	-1924671 when 5480,
	-1925324 when 5481,
	-1925977 when 5482,
	-1926628 when 5483,
	-1927278 when 5484,
	-1927927 when 5485,
	-1928574 when 5486,
	-1929221 when 5487,
	-1929866 when 5488,
	-1930510 when 5489,
	-1931153 when 5490,
	-1931795 when 5491,
	-1932435 when 5492,
	-1933074 when 5493,
	-1933712 when 5494,
	-1934349 when 5495,
	-1934985 when 5496,
	-1935619 when 5497,
	-1936253 when 5498,
	-1936885 when 5499,
	-1937516 when 5500,
	-1938146 when 5501,
	-1938774 when 5502,
	-1939401 when 5503,
	-1940028 when 5504,
	-1940652 when 5505,
	-1941276 when 5506,
	-1941899 when 5507,
	-1942520 when 5508,
	-1943140 when 5509,
	-1943759 when 5510,
	-1944377 when 5511,
	-1944993 when 5512,
	-1945609 when 5513,
	-1946223 when 5514,
	-1946836 when 5515,
	-1947448 when 5516,
	-1948058 when 5517,
	-1948668 when 5518,
	-1949276 when 5519,
	-1949883 when 5520,
	-1950488 when 5521,
	-1951093 when 5522,
	-1951696 when 5523,
	-1952298 when 5524,
	-1952899 when 5525,
	-1953499 when 5526,
	-1954097 when 5527,
	-1954695 when 5528,
	-1955291 when 5529,
	-1955886 when 5530,
	-1956479 when 5531,
	-1957072 when 5532,
	-1957663 when 5533,
	-1958253 when 5534,
	-1958842 when 5535,
	-1959430 when 5536,
	-1960016 when 5537,
	-1960601 when 5538,
	-1961186 when 5539,
	-1961768 when 5540,
	-1962350 when 5541,
	-1962930 when 5542,
	-1963509 when 5543,
	-1964087 when 5544,
	-1964664 when 5545,
	-1965240 when 5546,
	-1965814 when 5547,
	-1966387 when 5548,
	-1966959 when 5549,
	-1967530 when 5550,
	-1968099 when 5551,
	-1968668 when 5552,
	-1969235 when 5553,
	-1969800 when 5554,
	-1970365 when 5555,
	-1970929 when 5556,
	-1971491 when 5557,
	-1972052 when 5558,
	-1972611 when 5559,
	-1973170 when 5560,
	-1973727 when 5561,
	-1974283 when 5562,
	-1974838 when 5563,
	-1975392 when 5564,
	-1975944 when 5565,
	-1976496 when 5566,
	-1977046 when 5567,
	-1977594 when 5568,
	-1978142 when 5569,
	-1978688 when 5570,
	-1979234 when 5571,
	-1979777 when 5572,
	-1980320 when 5573,
	-1980862 when 5574,
	-1981402 when 5575,
	-1981941 when 5576,
	-1982479 when 5577,
	-1983015 when 5578,
	-1983551 when 5579,
	-1984085 when 5580,
	-1984618 when 5581,
	-1985149 when 5582,
	-1985680 when 5583,
	-1986209 when 5584,
	-1986737 when 5585,
	-1987264 when 5586,
	-1987789 when 5587,
	-1988314 when 5588,
	-1988837 when 5589,
	-1989359 when 5590,
	-1989879 when 5591,
	-1990399 when 5592,
	-1990917 when 5593,
	-1991434 when 5594,
	-1991950 when 5595,
	-1992464 when 5596,
	-1992978 when 5597,
	-1993490 when 5598,
	-1994000 when 5599,
	-1994510 when 5600,
	-1995018 when 5601,
	-1995526 when 5602,
	-1996031 when 5603,
	-1996536 when 5604,
	-1997040 when 5605,
	-1997542 when 5606,
	-1998043 when 5607,
	-1998543 when 5608,
	-1999041 when 5609,
	-1999538 when 5610,
	-2000034 when 5611,
	-2000529 when 5612,
	-2001023 when 5613,
	-2001515 when 5614,
	-2002006 when 5615,
	-2002496 when 5616,
	-2002985 when 5617,
	-2003472 when 5618,
	-2003958 when 5619,
	-2004443 when 5620,
	-2004927 when 5621,
	-2005409 when 5622,
	-2005891 when 5623,
	-2006371 when 5624,
	-2006849 when 5625,
	-2007327 when 5626,
	-2007803 when 5627,
	-2008278 when 5628,
	-2008752 when 5629,
	-2009224 when 5630,
	-2009696 when 5631,
	-2010166 when 5632,
	-2010635 when 5633,
	-2011102 when 5634,
	-2011569 when 5635,
	-2012034 when 5636,
	-2012498 when 5637,
	-2012960 when 5638,
	-2013422 when 5639,
	-2013882 when 5640,
	-2014341 when 5641,
	-2014798 when 5642,
	-2015255 when 5643,
	-2015710 when 5644,
	-2016164 when 5645,
	-2016617 when 5646,
	-2017068 when 5647,
	-2017518 when 5648,
	-2017967 when 5649,
	-2018415 when 5650,
	-2018861 when 5651,
	-2019307 when 5652,
	-2019751 when 5653,
	-2020193 when 5654,
	-2020635 when 5655,
	-2021075 when 5656,
	-2021514 when 5657,
	-2021952 when 5658,
	-2022388 when 5659,
	-2022824 when 5660,
	-2023258 when 5661,
	-2023690 when 5662,
	-2024122 when 5663,
	-2024552 when 5664,
	-2024981 when 5665,
	-2025409 when 5666,
	-2025835 when 5667,
	-2026261 when 5668,
	-2026685 when 5669,
	-2027107 when 5670,
	-2027529 when 5671,
	-2027949 when 5672,
	-2028368 when 5673,
	-2028786 when 5674,
	-2029202 when 5675,
	-2029618 when 5676,
	-2030032 when 5677,
	-2030444 when 5678,
	-2030856 when 5679,
	-2031266 when 5680,
	-2031675 when 5681,
	-2032083 when 5682,
	-2032489 when 5683,
	-2032895 when 5684,
	-2033299 when 5685,
	-2033701 when 5686,
	-2034103 when 5687,
	-2034503 when 5688,
	-2034902 when 5689,
	-2035300 when 5690,
	-2035696 when 5691,
	-2036091 when 5692,
	-2036485 when 5693,
	-2036878 when 5694,
	-2037269 when 5695,
	-2037659 when 5696,
	-2038048 when 5697,
	-2038436 when 5698,
	-2038822 when 5699,
	-2039208 when 5700,
	-2039591 when 5701,
	-2039974 when 5702,
	-2040355 when 5703,
	-2040735 when 5704,
	-2041114 when 5705,
	-2041492 when 5706,
	-2041868 when 5707,
	-2042243 when 5708,
	-2042617 when 5709,
	-2042990 when 5710,
	-2043361 when 5711,
	-2043731 when 5712,
	-2044100 when 5713,
	-2044467 when 5714,
	-2044833 when 5715,
	-2045198 when 5716,
	-2045562 when 5717,
	-2045925 when 5718,
	-2046286 when 5719,
	-2046646 when 5720,
	-2047004 when 5721,
	-2047362 when 5722,
	-2047718 when 5723,
	-2048073 when 5724,
	-2048427 when 5725,
	-2048779 when 5726,
	-2049130 when 5727,
	-2049480 when 5728,
	-2049828 when 5729,
	-2050176 when 5730,
	-2050522 when 5731,
	-2050866 when 5732,
	-2051210 when 5733,
	-2051552 when 5734,
	-2051893 when 5735,
	-2052233 when 5736,
	-2052571 when 5737,
	-2052909 when 5738,
	-2053244 when 5739,
	-2053579 when 5740,
	-2053912 when 5741,
	-2054245 when 5742,
	-2054575 when 5743,
	-2054905 when 5744,
	-2055233 when 5745,
	-2055560 when 5746,
	-2055886 when 5747,
	-2056211 when 5748,
	-2056534 when 5749,
	-2056856 when 5750,
	-2057177 when 5751,
	-2057496 when 5752,
	-2057814 when 5753,
	-2058131 when 5754,
	-2058447 when 5755,
	-2058761 when 5756,
	-2059074 when 5757,
	-2059386 when 5758,
	-2059696 when 5759,
	-2060006 when 5760,
	-2060314 when 5761,
	-2060620 when 5762,
	-2060926 when 5763,
	-2061230 when 5764,
	-2061533 when 5765,
	-2061835 when 5766,
	-2062135 when 5767,
	-2062434 when 5768,
	-2062732 when 5769,
	-2063028 when 5770,
	-2063324 when 5771,
	-2063618 when 5772,
	-2063910 when 5773,
	-2064202 when 5774,
	-2064492 when 5775,
	-2064781 when 5776,
	-2065069 when 5777,
	-2065355 when 5778,
	-2065640 when 5779,
	-2065924 when 5780,
	-2066207 when 5781,
	-2066488 when 5782,
	-2066768 when 5783,
	-2067047 when 5784,
	-2067324 when 5785,
	-2067600 when 5786,
	-2067875 when 5787,
	-2068149 when 5788,
	-2068421 when 5789,
	-2068692 when 5790,
	-2068962 when 5791,
	-2069230 when 5792,
	-2069498 when 5793,
	-2069764 when 5794,
	-2070028 when 5795,
	-2070292 when 5796,
	-2070554 when 5797,
	-2070815 when 5798,
	-2071074 when 5799,
	-2071333 when 5800,
	-2071590 when 5801,
	-2071845 when 5802,
	-2072100 when 5803,
	-2072353 when 5804,
	-2072605 when 5805,
	-2072856 when 5806,
	-2073105 when 5807,
	-2073353 when 5808,
	-2073600 when 5809,
	-2073845 when 5810,
	-2074090 when 5811,
	-2074332 when 5812,
	-2074574 when 5813,
	-2074815 when 5814,
	-2075054 when 5815,
	-2075292 when 5816,
	-2075528 when 5817,
	-2075763 when 5818,
	-2075997 when 5819,
	-2076230 when 5820,
	-2076462 when 5821,
	-2076692 when 5822,
	-2076921 when 5823,
	-2077148 when 5824,
	-2077374 when 5825,
	-2077600 when 5826,
	-2077823 when 5827,
	-2078046 when 5828,
	-2078267 when 5829,
	-2078487 when 5830,
	-2078705 when 5831,
	-2078923 when 5832,
	-2079139 when 5833,
	-2079354 when 5834,
	-2079567 when 5835,
	-2079779 when 5836,
	-2079990 when 5837,
	-2080200 when 5838,
	-2080408 when 5839,
	-2080615 when 5840,
	-2080821 when 5841,
	-2081026 when 5842,
	-2081229 when 5843,
	-2081431 when 5844,
	-2081631 when 5845,
	-2081831 when 5846,
	-2082029 when 5847,
	-2082226 when 5848,
	-2082421 when 5849,
	-2082616 when 5850,
	-2082808 when 5851,
	-2083000 when 5852,
	-2083191 when 5853,
	-2083380 when 5854,
	-2083567 when 5855,
	-2083754 when 5856,
	-2083939 when 5857,
	-2084123 when 5858,
	-2084306 when 5859,
	-2084487 when 5860,
	-2084667 when 5861,
	-2084846 when 5862,
	-2085024 when 5863,
	-2085200 when 5864,
	-2085375 when 5865,
	-2085549 when 5866,
	-2085721 when 5867,
	-2085892 when 5868,
	-2086062 when 5869,
	-2086230 when 5870,
	-2086398 when 5871,
	-2086564 when 5872,
	-2086728 when 5873,
	-2086892 when 5874,
	-2087054 when 5875,
	-2087214 when 5876,
	-2087374 when 5877,
	-2087532 when 5878,
	-2087689 when 5879,
	-2087845 when 5880,
	-2087999 when 5881,
	-2088152 when 5882,
	-2088304 when 5883,
	-2088454 when 5884,
	-2088604 when 5885,
	-2088752 when 5886,
	-2088898 when 5887,
	-2089044 when 5888,
	-2089188 when 5889,
	-2089330 when 5890,
	-2089472 when 5891,
	-2089612 when 5892,
	-2089751 when 5893,
	-2089889 when 5894,
	-2090025 when 5895,
	-2090160 when 5896,
	-2090294 when 5897,
	-2090426 when 5898,
	-2090557 when 5899,
	-2090687 when 5900,
	-2090816 when 5901,
	-2090943 when 5902,
	-2091069 when 5903,
	-2091194 when 5904,
	-2091317 when 5905,
	-2091439 when 5906,
	-2091560 when 5907,
	-2091680 when 5908,
	-2091798 when 5909,
	-2091915 when 5910,
	-2092031 when 5911,
	-2092145 when 5912,
	-2092258 when 5913,
	-2092370 when 5914,
	-2092481 when 5915,
	-2092590 when 5916,
	-2092698 when 5917,
	-2092804 when 5918,
	-2092910 when 5919,
	-2093014 when 5920,
	-2093117 when 5921,
	-2093218 when 5922,
	-2093318 when 5923,
	-2093417 when 5924,
	-2093515 when 5925,
	-2093611 when 5926,
	-2093706 when 5927,
	-2093800 when 5928,
	-2093892 when 5929,
	-2093983 when 5930,
	-2094073 when 5931,
	-2094162 when 5932,
	-2094249 when 5933,
	-2094335 when 5934,
	-2094420 when 5935,
	-2094503 when 5936,
	-2094585 when 5937,
	-2094666 when 5938,
	-2094746 when 5939,
	-2094824 when 5940,
	-2094901 when 5941,
	-2094976 when 5942,
	-2095051 when 5943,
	-2095124 when 5944,
	-2095196 when 5945,
	-2095266 when 5946,
	-2095335 when 5947,
	-2095403 when 5948,
	-2095470 when 5949,
	-2095535 when 5950,
	-2095599 when 5951,
	-2095662 when 5952,
	-2095723 when 5953,
	-2095783 when 5954,
	-2095842 when 5955,
	-2095900 when 5956,
	-2095956 when 5957,
	-2096011 when 5958,
	-2096065 when 5959,
	-2096117 when 5960,
	-2096168 when 5961,
	-2096218 when 5962,
	-2096267 when 5963,
	-2096314 when 5964,
	-2096360 when 5965,
	-2096404 when 5966,
	-2096448 when 5967,
	-2096490 when 5968,
	-2096530 when 5969,
	-2096570 when 5970,
	-2096608 when 5971,
	-2096645 when 5972,
	-2096680 when 5973,
	-2096715 when 5974,
	-2096748 when 5975,
	-2096779 when 5976,
	-2096810 when 5977,
	-2096839 when 5978,
	-2096867 when 5979,
	-2096893 when 5980,
	-2096919 when 5981,
	-2096942 when 5982,
	-2096965 when 5983,
	-2096986 when 5984,
	-2097006 when 5985,
	-2097025 when 5986,
	-2097043 when 5987,
	-2097059 when 5988,
	-2097074 when 5989,
	-2097087 when 5990,
	-2097100 when 5991,
	-2097111 when 5992,
	-2097120 when 5993,
	-2097129 when 5994,
	-2097136 when 5995,
	-2097142 when 5996,
	-2097146 when 5997,
	-2097149 when 5998,
	-2097151 when 5999,
	-2097152 when 6000,
	-2097151 when 6001,
	-2097149 when 6002,
	-2097146 when 6003,
	-2097142 when 6004,
	-2097136 when 6005,
	-2097129 when 6006,
	-2097120 when 6007,
	-2097111 when 6008,
	-2097100 when 6009,
	-2097087 when 6010,
	-2097074 when 6011,
	-2097059 when 6012,
	-2097043 when 6013,
	-2097025 when 6014,
	-2097006 when 6015,
	-2096986 when 6016,
	-2096965 when 6017,
	-2096942 when 6018,
	-2096919 when 6019,
	-2096893 when 6020,
	-2096867 when 6021,
	-2096839 when 6022,
	-2096810 when 6023,
	-2096779 when 6024,
	-2096748 when 6025,
	-2096715 when 6026,
	-2096680 when 6027,
	-2096645 when 6028,
	-2096608 when 6029,
	-2096570 when 6030,
	-2096530 when 6031,
	-2096490 when 6032,
	-2096448 when 6033,
	-2096404 when 6034,
	-2096360 when 6035,
	-2096314 when 6036,
	-2096267 when 6037,
	-2096218 when 6038,
	-2096168 when 6039,
	-2096117 when 6040,
	-2096065 when 6041,
	-2096011 when 6042,
	-2095956 when 6043,
	-2095900 when 6044,
	-2095842 when 6045,
	-2095783 when 6046,
	-2095723 when 6047,
	-2095662 when 6048,
	-2095599 when 6049,
	-2095535 when 6050,
	-2095470 when 6051,
	-2095403 when 6052,
	-2095335 when 6053,
	-2095266 when 6054,
	-2095196 when 6055,
	-2095124 when 6056,
	-2095051 when 6057,
	-2094976 when 6058,
	-2094901 when 6059,
	-2094824 when 6060,
	-2094746 when 6061,
	-2094666 when 6062,
	-2094585 when 6063,
	-2094503 when 6064,
	-2094420 when 6065,
	-2094335 when 6066,
	-2094249 when 6067,
	-2094162 when 6068,
	-2094073 when 6069,
	-2093983 when 6070,
	-2093892 when 6071,
	-2093800 when 6072,
	-2093706 when 6073,
	-2093611 when 6074,
	-2093515 when 6075,
	-2093417 when 6076,
	-2093318 when 6077,
	-2093218 when 6078,
	-2093117 when 6079,
	-2093014 when 6080,
	-2092910 when 6081,
	-2092804 when 6082,
	-2092698 when 6083,
	-2092590 when 6084,
	-2092481 when 6085,
	-2092370 when 6086,
	-2092258 when 6087,
	-2092145 when 6088,
	-2092031 when 6089,
	-2091915 when 6090,
	-2091798 when 6091,
	-2091680 when 6092,
	-2091560 when 6093,
	-2091439 when 6094,
	-2091317 when 6095,
	-2091194 when 6096,
	-2091069 when 6097,
	-2090943 when 6098,
	-2090816 when 6099,
	-2090687 when 6100,
	-2090557 when 6101,
	-2090426 when 6102,
	-2090294 when 6103,
	-2090160 when 6104,
	-2090025 when 6105,
	-2089889 when 6106,
	-2089751 when 6107,
	-2089612 when 6108,
	-2089472 when 6109,
	-2089330 when 6110,
	-2089188 when 6111,
	-2089044 when 6112,
	-2088898 when 6113,
	-2088752 when 6114,
	-2088604 when 6115,
	-2088454 when 6116,
	-2088304 when 6117,
	-2088152 when 6118,
	-2087999 when 6119,
	-2087845 when 6120,
	-2087689 when 6121,
	-2087532 when 6122,
	-2087374 when 6123,
	-2087214 when 6124,
	-2087054 when 6125,
	-2086892 when 6126,
	-2086728 when 6127,
	-2086564 when 6128,
	-2086398 when 6129,
	-2086230 when 6130,
	-2086062 when 6131,
	-2085892 when 6132,
	-2085721 when 6133,
	-2085549 when 6134,
	-2085375 when 6135,
	-2085200 when 6136,
	-2085024 when 6137,
	-2084846 when 6138,
	-2084667 when 6139,
	-2084487 when 6140,
	-2084306 when 6141,
	-2084123 when 6142,
	-2083939 when 6143,
	-2083754 when 6144,
	-2083567 when 6145,
	-2083380 when 6146,
	-2083191 when 6147,
	-2083000 when 6148,
	-2082808 when 6149,
	-2082616 when 6150,
	-2082421 when 6151,
	-2082226 when 6152,
	-2082029 when 6153,
	-2081831 when 6154,
	-2081631 when 6155,
	-2081431 when 6156,
	-2081229 when 6157,
	-2081026 when 6158,
	-2080821 when 6159,
	-2080615 when 6160,
	-2080408 when 6161,
	-2080200 when 6162,
	-2079990 when 6163,
	-2079779 when 6164,
	-2079567 when 6165,
	-2079354 when 6166,
	-2079139 when 6167,
	-2078923 when 6168,
	-2078705 when 6169,
	-2078487 when 6170,
	-2078267 when 6171,
	-2078046 when 6172,
	-2077823 when 6173,
	-2077600 when 6174,
	-2077374 when 6175,
	-2077148 when 6176,
	-2076921 when 6177,
	-2076692 when 6178,
	-2076462 when 6179,
	-2076230 when 6180,
	-2075997 when 6181,
	-2075763 when 6182,
	-2075528 when 6183,
	-2075292 when 6184,
	-2075054 when 6185,
	-2074815 when 6186,
	-2074574 when 6187,
	-2074332 when 6188,
	-2074090 when 6189,
	-2073845 when 6190,
	-2073600 when 6191,
	-2073353 when 6192,
	-2073105 when 6193,
	-2072856 when 6194,
	-2072605 when 6195,
	-2072353 when 6196,
	-2072100 when 6197,
	-2071845 when 6198,
	-2071590 when 6199,
	-2071333 when 6200,
	-2071074 when 6201,
	-2070815 when 6202,
	-2070554 when 6203,
	-2070292 when 6204,
	-2070028 when 6205,
	-2069764 when 6206,
	-2069498 when 6207,
	-2069230 when 6208,
	-2068962 when 6209,
	-2068692 when 6210,
	-2068421 when 6211,
	-2068149 when 6212,
	-2067875 when 6213,
	-2067600 when 6214,
	-2067324 when 6215,
	-2067047 when 6216,
	-2066768 when 6217,
	-2066488 when 6218,
	-2066207 when 6219,
	-2065924 when 6220,
	-2065640 when 6221,
	-2065355 when 6222,
	-2065069 when 6223,
	-2064781 when 6224,
	-2064492 when 6225,
	-2064202 when 6226,
	-2063910 when 6227,
	-2063618 when 6228,
	-2063324 when 6229,
	-2063028 when 6230,
	-2062732 when 6231,
	-2062434 when 6232,
	-2062135 when 6233,
	-2061835 when 6234,
	-2061533 when 6235,
	-2061230 when 6236,
	-2060926 when 6237,
	-2060620 when 6238,
	-2060314 when 6239,
	-2060006 when 6240,
	-2059696 when 6241,
	-2059386 when 6242,
	-2059074 when 6243,
	-2058761 when 6244,
	-2058447 when 6245,
	-2058131 when 6246,
	-2057814 when 6247,
	-2057496 when 6248,
	-2057177 when 6249,
	-2056856 when 6250,
	-2056534 when 6251,
	-2056211 when 6252,
	-2055886 when 6253,
	-2055560 when 6254,
	-2055233 when 6255,
	-2054905 when 6256,
	-2054575 when 6257,
	-2054245 when 6258,
	-2053912 when 6259,
	-2053579 when 6260,
	-2053244 when 6261,
	-2052909 when 6262,
	-2052571 when 6263,
	-2052233 when 6264,
	-2051893 when 6265,
	-2051552 when 6266,
	-2051210 when 6267,
	-2050866 when 6268,
	-2050522 when 6269,
	-2050176 when 6270,
	-2049828 when 6271,
	-2049480 when 6272,
	-2049130 when 6273,
	-2048779 when 6274,
	-2048427 when 6275,
	-2048073 when 6276,
	-2047718 when 6277,
	-2047362 when 6278,
	-2047004 when 6279,
	-2046646 when 6280,
	-2046286 when 6281,
	-2045925 when 6282,
	-2045562 when 6283,
	-2045198 when 6284,
	-2044833 when 6285,
	-2044467 when 6286,
	-2044100 when 6287,
	-2043731 when 6288,
	-2043361 when 6289,
	-2042990 when 6290,
	-2042617 when 6291,
	-2042243 when 6292,
	-2041868 when 6293,
	-2041492 when 6294,
	-2041114 when 6295,
	-2040735 when 6296,
	-2040355 when 6297,
	-2039974 when 6298,
	-2039591 when 6299,
	-2039208 when 6300,
	-2038822 when 6301,
	-2038436 when 6302,
	-2038048 when 6303,
	-2037659 when 6304,
	-2037269 when 6305,
	-2036878 when 6306,
	-2036485 when 6307,
	-2036091 when 6308,
	-2035696 when 6309,
	-2035300 when 6310,
	-2034902 when 6311,
	-2034503 when 6312,
	-2034103 when 6313,
	-2033701 when 6314,
	-2033299 when 6315,
	-2032895 when 6316,
	-2032489 when 6317,
	-2032083 when 6318,
	-2031675 when 6319,
	-2031266 when 6320,
	-2030856 when 6321,
	-2030444 when 6322,
	-2030032 when 6323,
	-2029618 when 6324,
	-2029202 when 6325,
	-2028786 when 6326,
	-2028368 when 6327,
	-2027949 when 6328,
	-2027529 when 6329,
	-2027107 when 6330,
	-2026685 when 6331,
	-2026261 when 6332,
	-2025835 when 6333,
	-2025409 when 6334,
	-2024981 when 6335,
	-2024552 when 6336,
	-2024122 when 6337,
	-2023690 when 6338,
	-2023258 when 6339,
	-2022824 when 6340,
	-2022388 when 6341,
	-2021952 when 6342,
	-2021514 when 6343,
	-2021075 when 6344,
	-2020635 when 6345,
	-2020193 when 6346,
	-2019751 when 6347,
	-2019307 when 6348,
	-2018861 when 6349,
	-2018415 when 6350,
	-2017967 when 6351,
	-2017518 when 6352,
	-2017068 when 6353,
	-2016617 when 6354,
	-2016164 when 6355,
	-2015710 when 6356,
	-2015255 when 6357,
	-2014798 when 6358,
	-2014341 when 6359,
	-2013882 when 6360,
	-2013422 when 6361,
	-2012960 when 6362,
	-2012498 when 6363,
	-2012034 when 6364,
	-2011569 when 6365,
	-2011102 when 6366,
	-2010635 when 6367,
	-2010166 when 6368,
	-2009696 when 6369,
	-2009224 when 6370,
	-2008752 when 6371,
	-2008278 when 6372,
	-2007803 when 6373,
	-2007327 when 6374,
	-2006849 when 6375,
	-2006371 when 6376,
	-2005891 when 6377,
	-2005409 when 6378,
	-2004927 when 6379,
	-2004443 when 6380,
	-2003958 when 6381,
	-2003472 when 6382,
	-2002985 when 6383,
	-2002496 when 6384,
	-2002006 when 6385,
	-2001515 when 6386,
	-2001023 when 6387,
	-2000529 when 6388,
	-2000034 when 6389,
	-1999538 when 6390,
	-1999041 when 6391,
	-1998543 when 6392,
	-1998043 when 6393,
	-1997542 when 6394,
	-1997040 when 6395,
	-1996536 when 6396,
	-1996031 when 6397,
	-1995526 when 6398,
	-1995018 when 6399,
	-1994510 when 6400,
	-1994000 when 6401,
	-1993490 when 6402,
	-1992978 when 6403,
	-1992464 when 6404,
	-1991950 when 6405,
	-1991434 when 6406,
	-1990917 when 6407,
	-1990399 when 6408,
	-1989879 when 6409,
	-1989359 when 6410,
	-1988837 when 6411,
	-1988314 when 6412,
	-1987789 when 6413,
	-1987264 when 6414,
	-1986737 when 6415,
	-1986209 when 6416,
	-1985680 when 6417,
	-1985149 when 6418,
	-1984618 when 6419,
	-1984085 when 6420,
	-1983551 when 6421,
	-1983015 when 6422,
	-1982479 when 6423,
	-1981941 when 6424,
	-1981402 when 6425,
	-1980862 when 6426,
	-1980320 when 6427,
	-1979777 when 6428,
	-1979234 when 6429,
	-1978688 when 6430,
	-1978142 when 6431,
	-1977594 when 6432,
	-1977046 when 6433,
	-1976496 when 6434,
	-1975944 when 6435,
	-1975392 when 6436,
	-1974838 when 6437,
	-1974283 when 6438,
	-1973727 when 6439,
	-1973170 when 6440,
	-1972611 when 6441,
	-1972052 when 6442,
	-1971491 when 6443,
	-1970929 when 6444,
	-1970365 when 6445,
	-1969800 when 6446,
	-1969235 when 6447,
	-1968668 when 6448,
	-1968099 when 6449,
	-1967530 when 6450,
	-1966959 when 6451,
	-1966387 when 6452,
	-1965814 when 6453,
	-1965240 when 6454,
	-1964664 when 6455,
	-1964087 when 6456,
	-1963509 when 6457,
	-1962930 when 6458,
	-1962350 when 6459,
	-1961768 when 6460,
	-1961186 when 6461,
	-1960601 when 6462,
	-1960016 when 6463,
	-1959430 when 6464,
	-1958842 when 6465,
	-1958253 when 6466,
	-1957663 when 6467,
	-1957072 when 6468,
	-1956479 when 6469,
	-1955886 when 6470,
	-1955291 when 6471,
	-1954695 when 6472,
	-1954097 when 6473,
	-1953499 when 6474,
	-1952899 when 6475,
	-1952298 when 6476,
	-1951696 when 6477,
	-1951093 when 6478,
	-1950488 when 6479,
	-1949883 when 6480,
	-1949276 when 6481,
	-1948668 when 6482,
	-1948058 when 6483,
	-1947448 when 6484,
	-1946836 when 6485,
	-1946223 when 6486,
	-1945609 when 6487,
	-1944993 when 6488,
	-1944377 when 6489,
	-1943759 when 6490,
	-1943140 when 6491,
	-1942520 when 6492,
	-1941899 when 6493,
	-1941276 when 6494,
	-1940652 when 6495,
	-1940028 when 6496,
	-1939401 when 6497,
	-1938774 when 6498,
	-1938146 when 6499,
	-1937516 when 6500,
	-1936885 when 6501,
	-1936253 when 6502,
	-1935619 when 6503,
	-1934985 when 6504,
	-1934349 when 6505,
	-1933712 when 6506,
	-1933074 when 6507,
	-1932435 when 6508,
	-1931795 when 6509,
	-1931153 when 6510,
	-1930510 when 6511,
	-1929866 when 6512,
	-1929221 when 6513,
	-1928574 when 6514,
	-1927927 when 6515,
	-1927278 when 6516,
	-1926628 when 6517,
	-1925977 when 6518,
	-1925324 when 6519,
	-1924671 when 6520,
	-1924016 when 6521,
	-1923360 when 6522,
	-1922703 when 6523,
	-1922045 when 6524,
	-1921385 when 6525,
	-1920725 when 6526,
	-1920063 when 6527,
	-1919400 when 6528,
	-1918736 when 6529,
	-1918070 when 6530,
	-1917404 when 6531,
	-1916736 when 6532,
	-1916067 when 6533,
	-1915397 when 6534,
	-1914725 when 6535,
	-1914053 when 6536,
	-1913379 when 6537,
	-1912704 when 6538,
	-1912028 when 6539,
	-1911351 when 6540,
	-1910673 when 6541,
	-1909993 when 6542,
	-1909312 when 6543,
	-1908631 when 6544,
	-1907947 when 6545,
	-1907263 when 6546,
	-1906578 when 6547,
	-1905891 when 6548,
	-1905203 when 6549,
	-1904514 when 6550,
	-1903824 when 6551,
	-1903133 when 6552,
	-1902440 when 6553,
	-1901747 when 6554,
	-1901052 when 6555,
	-1900356 when 6556,
	-1899658 when 6557,
	-1898960 when 6558,
	-1898261 when 6559,
	-1897560 when 6560,
	-1896858 when 6561,
	-1896155 when 6562,
	-1895451 when 6563,
	-1894745 when 6564,
	-1894039 when 6565,
	-1893331 when 6566,
	-1892622 when 6567,
	-1891912 when 6568,
	-1891201 when 6569,
	-1890488 when 6570,
	-1889775 when 6571,
	-1889060 when 6572,
	-1888344 when 6573,
	-1887627 when 6574,
	-1886909 when 6575,
	-1886190 when 6576,
	-1885469 when 6577,
	-1884747 when 6578,
	-1884024 when 6579,
	-1883300 when 6580,
	-1882575 when 6581,
	-1881849 when 6582,
	-1881121 when 6583,
	-1880393 when 6584,
	-1879663 when 6585,
	-1878932 when 6586,
	-1878200 when 6587,
	-1877466 when 6588,
	-1876732 when 6589,
	-1875996 when 6590,
	-1875259 when 6591,
	-1874521 when 6592,
	-1873782 when 6593,
	-1873042 when 6594,
	-1872301 when 6595,
	-1871558 when 6596,
	-1870814 when 6597,
	-1870069 when 6598,
	-1869323 when 6599,
	-1868576 when 6600,
	-1867828 when 6601,
	-1867078 when 6602,
	-1866328 when 6603,
	-1865576 when 6604,
	-1864823 when 6605,
	-1864069 when 6606,
	-1863314 when 6607,
	-1862557 when 6608,
	-1861800 when 6609,
	-1861041 when 6610,
	-1860281 when 6611,
	-1859520 when 6612,
	-1858758 when 6613,
	-1857995 when 6614,
	-1857230 when 6615,
	-1856465 when 6616,
	-1855698 when 6617,
	-1854930 when 6618,
	-1854161 when 6619,
	-1853391 when 6620,
	-1852620 when 6621,
	-1851847 when 6622,
	-1851074 when 6623,
	-1850299 when 6624,
	-1849523 when 6625,
	-1848746 when 6626,
	-1847968 when 6627,
	-1847188 when 6628,
	-1846408 when 6629,
	-1845627 when 6630,
	-1844844 when 6631,
	-1844060 when 6632,
	-1843275 when 6633,
	-1842489 when 6634,
	-1841702 when 6635,
	-1840913 when 6636,
	-1840124 when 6637,
	-1839333 when 6638,
	-1838541 when 6639,
	-1837748 when 6640,
	-1836954 when 6641,
	-1836159 when 6642,
	-1835363 when 6643,
	-1834565 when 6644,
	-1833767 when 6645,
	-1832967 when 6646,
	-1832166 when 6647,
	-1831364 when 6648,
	-1830561 when 6649,
	-1829757 when 6650,
	-1828951 when 6651,
	-1828145 when 6652,
	-1827337 when 6653,
	-1826528 when 6654,
	-1825719 when 6655,
	-1824908 when 6656,
	-1824095 when 6657,
	-1823282 when 6658,
	-1822468 when 6659,
	-1821652 when 6660,
	-1820836 when 6661,
	-1820018 when 6662,
	-1819199 when 6663,
	-1818379 when 6664,
	-1817558 when 6665,
	-1816736 when 6666,
	-1815912 when 6667,
	-1815088 when 6668,
	-1814262 when 6669,
	-1813436 when 6670,
	-1812608 when 6671,
	-1811779 when 6672,
	-1810949 when 6673,
	-1810117 when 6674,
	-1809285 when 6675,
	-1808452 when 6676,
	-1807617 when 6677,
	-1806782 when 6678,
	-1805945 when 6679,
	-1805107 when 6680,
	-1804268 when 6681,
	-1803428 when 6682,
	-1802587 when 6683,
	-1801744 when 6684,
	-1800901 when 6685,
	-1800056 when 6686,
	-1799211 when 6687,
	-1798364 when 6688,
	-1797516 when 6689,
	-1796667 when 6690,
	-1795817 when 6691,
	-1794966 when 6692,
	-1794113 when 6693,
	-1793260 when 6694,
	-1792405 when 6695,
	-1791550 when 6696,
	-1790693 when 6697,
	-1789835 when 6698,
	-1788976 when 6699,
	-1788116 when 6700,
	-1787255 when 6701,
	-1786393 when 6702,
	-1785529 when 6703,
	-1784665 when 6704,
	-1783799 when 6705,
	-1782933 when 6706,
	-1782065 when 6707,
	-1781196 when 6708,
	-1780326 when 6709,
	-1779455 when 6710,
	-1778583 when 6711,
	-1777709 when 6712,
	-1776835 when 6713,
	-1775960 when 6714,
	-1775083 when 6715,
	-1774205 when 6716,
	-1773327 when 6717,
	-1772447 when 6718,
	-1771566 when 6719,
	-1770684 when 6720,
	-1769801 when 6721,
	-1768917 when 6722,
	-1768031 when 6723,
	-1767145 when 6724,
	-1766258 when 6725,
	-1765369 when 6726,
	-1764479 when 6727,
	-1763589 when 6728,
	-1762697 when 6729,
	-1761804 when 6730,
	-1760910 when 6731,
	-1760015 when 6732,
	-1759119 when 6733,
	-1758221 when 6734,
	-1757323 when 6735,
	-1756424 when 6736,
	-1755523 when 6737,
	-1754622 when 6738,
	-1753719 when 6739,
	-1752815 when 6740,
	-1751910 when 6741,
	-1751004 when 6742,
	-1750097 when 6743,
	-1749189 when 6744,
	-1748280 when 6745,
	-1747370 when 6746,
	-1746459 when 6747,
	-1745546 when 6748,
	-1744633 when 6749,
	-1743718 when 6750,
	-1742803 when 6751,
	-1741886 when 6752,
	-1740968 when 6753,
	-1740049 when 6754,
	-1739129 when 6755,
	-1738208 when 6756,
	-1737286 when 6757,
	-1736363 when 6758,
	-1735439 when 6759,
	-1734514 when 6760,
	-1733587 when 6761,
	-1732660 when 6762,
	-1731731 when 6763,
	-1730802 when 6764,
	-1729871 when 6765,
	-1728940 when 6766,
	-1728007 when 6767,
	-1727073 when 6768,
	-1726138 when 6769,
	-1725202 when 6770,
	-1724265 when 6771,
	-1723327 when 6772,
	-1722388 when 6773,
	-1721448 when 6774,
	-1720507 when 6775,
	-1719564 when 6776,
	-1718621 when 6777,
	-1717676 when 6778,
	-1716731 when 6779,
	-1715784 when 6780,
	-1714837 when 6781,
	-1713888 when 6782,
	-1712938 when 6783,
	-1711987 when 6784,
	-1711036 when 6785,
	-1710083 when 6786,
	-1709129 when 6787,
	-1708174 when 6788,
	-1707218 when 6789,
	-1706261 when 6790,
	-1705302 when 6791,
	-1704343 when 6792,
	-1703383 when 6793,
	-1702422 when 6794,
	-1701459 when 6795,
	-1700496 when 6796,
	-1699531 when 6797,
	-1698566 when 6798,
	-1697599 when 6799,
	-1696632 when 6800,
	-1695663 when 6801,
	-1694693 when 6802,
	-1693722 when 6803,
	-1692751 when 6804,
	-1691778 when 6805,
	-1690804 when 6806,
	-1689829 when 6807,
	-1688853 when 6808,
	-1687876 when 6809,
	-1686898 when 6810,
	-1685919 when 6811,
	-1684939 when 6812,
	-1683958 when 6813,
	-1682975 when 6814,
	-1681992 when 6815,
	-1681008 when 6816,
	-1680022 when 6817,
	-1679036 when 6818,
	-1678049 when 6819,
	-1677060 when 6820,
	-1676071 when 6821,
	-1675080 when 6822,
	-1674089 when 6823,
	-1673096 when 6824,
	-1672103 when 6825,
	-1671108 when 6826,
	-1670112 when 6827,
	-1669116 when 6828,
	-1668118 when 6829,
	-1667119 when 6830,
	-1666119 when 6831,
	-1665119 when 6832,
	-1664117 when 6833,
	-1663114 when 6834,
	-1662110 when 6835,
	-1661105 when 6836,
	-1660099 when 6837,
	-1659092 when 6838,
	-1658084 when 6839,
	-1657075 when 6840,
	-1656065 when 6841,
	-1655054 when 6842,
	-1654042 when 6843,
	-1653029 when 6844,
	-1652015 when 6845,
	-1651000 when 6846,
	-1649984 when 6847,
	-1648966 when 6848,
	-1647948 when 6849,
	-1646929 when 6850,
	-1645909 when 6851,
	-1644888 when 6852,
	-1643865 when 6853,
	-1642842 when 6854,
	-1641818 when 6855,
	-1640792 when 6856,
	-1639766 when 6857,
	-1638739 when 6858,
	-1637711 when 6859,
	-1636681 when 6860,
	-1635651 when 6861,
	-1634619 when 6862,
	-1633587 when 6863,
	-1632554 when 6864,
	-1631519 when 6865,
	-1630484 when 6866,
	-1629448 when 6867,
	-1628410 when 6868,
	-1627372 when 6869,
	-1626332 when 6870,
	-1625292 when 6871,
	-1624251 when 6872,
	-1623208 when 6873,
	-1622165 when 6874,
	-1621120 when 6875,
	-1620075 when 6876,
	-1619029 when 6877,
	-1617981 when 6878,
	-1616933 when 6879,
	-1615883 when 6880,
	-1614833 when 6881,
	-1613782 when 6882,
	-1612729 when 6883,
	-1611676 when 6884,
	-1610621 when 6885,
	-1609566 when 6886,
	-1608510 when 6887,
	-1607452 when 6888,
	-1606394 when 6889,
	-1605335 when 6890,
	-1604274 when 6891,
	-1603213 when 6892,
	-1602151 when 6893,
	-1601087 when 6894,
	-1600023 when 6895,
	-1598958 when 6896,
	-1597892 when 6897,
	-1596824 when 6898,
	-1595756 when 6899,
	-1594687 when 6900,
	-1593617 when 6901,
	-1592546 when 6902,
	-1591473 when 6903,
	-1590400 when 6904,
	-1589326 when 6905,
	-1588251 when 6906,
	-1587175 when 6907,
	-1586098 when 6908,
	-1585020 when 6909,
	-1583941 when 6910,
	-1582861 when 6911,
	-1581780 when 6912,
	-1580698 when 6913,
	-1579615 when 6914,
	-1578531 when 6915,
	-1577446 when 6916,
	-1576360 when 6917,
	-1575273 when 6918,
	-1574186 when 6919,
	-1573097 when 6920,
	-1572007 when 6921,
	-1570916 when 6922,
	-1569825 when 6923,
	-1568732 when 6924,
	-1567639 when 6925,
	-1566544 when 6926,
	-1565448 when 6927,
	-1564352 when 6928,
	-1563254 when 6929,
	-1562156 when 6930,
	-1561057 when 6931,
	-1559956 when 6932,
	-1558855 when 6933,
	-1557753 when 6934,
	-1556649 when 6935,
	-1555545 when 6936,
	-1554440 when 6937,
	-1553334 when 6938,
	-1552227 when 6939,
	-1551119 when 6940,
	-1550010 when 6941,
	-1548900 when 6942,
	-1547789 when 6943,
	-1546677 when 6944,
	-1545564 when 6945,
	-1544451 when 6946,
	-1543336 when 6947,
	-1542220 when 6948,
	-1541103 when 6949,
	-1539986 when 6950,
	-1538867 when 6951,
	-1537748 when 6952,
	-1536627 when 6953,
	-1535506 when 6954,
	-1534384 when 6955,
	-1533261 when 6956,
	-1532136 when 6957,
	-1531011 when 6958,
	-1529885 when 6959,
	-1528758 when 6960,
	-1527630 when 6961,
	-1526501 when 6962,
	-1525371 when 6963,
	-1524240 when 6964,
	-1523109 when 6965,
	-1521976 when 6966,
	-1520842 when 6967,
	-1519708 when 6968,
	-1518572 when 6969,
	-1517436 when 6970,
	-1516298 when 6971,
	-1515160 when 6972,
	-1514021 when 6973,
	-1512881 when 6974,
	-1511740 when 6975,
	-1510598 when 6976,
	-1509455 when 6977,
	-1508311 when 6978,
	-1507166 when 6979,
	-1506020 when 6980,
	-1504873 when 6981,
	-1503726 when 6982,
	-1502577 when 6983,
	-1501428 when 6984,
	-1500277 when 6985,
	-1499126 when 6986,
	-1497974 when 6987,
	-1496820 when 6988,
	-1495666 when 6989,
	-1494511 when 6990,
	-1493355 when 6991,
	-1492198 when 6992,
	-1491041 when 6993,
	-1489882 when 6994,
	-1488722 when 6995,
	-1487562 when 6996,
	-1486400 when 6997,
	-1485238 when 6998,
	-1484075 when 6999,
	-1482910 when 7000,
	-1481745 when 7001,
	-1480579 when 7002,
	-1479412 when 7003,
	-1478244 when 7004,
	-1477076 when 7005,
	-1475906 when 7006,
	-1474735 when 7007,
	-1473564 when 7008,
	-1472391 when 7009,
	-1471218 when 7010,
	-1470044 when 7011,
	-1468869 when 7012,
	-1467693 when 7013,
	-1466516 when 7014,
	-1465338 when 7015,
	-1464159 when 7016,
	-1462979 when 7017,
	-1461799 when 7018,
	-1460617 when 7019,
	-1459435 when 7020,
	-1458252 when 7021,
	-1457067 when 7022,
	-1455882 when 7023,
	-1454696 when 7024,
	-1453510 when 7025,
	-1452322 when 7026,
	-1451133 when 7027,
	-1449944 when 7028,
	-1448753 when 7029,
	-1447562 when 7030,
	-1446370 when 7031,
	-1445176 when 7032,
	-1443982 when 7033,
	-1442787 when 7034,
	-1441592 when 7035,
	-1440395 when 7036,
	-1439197 when 7037,
	-1437999 when 7038,
	-1436800 when 7039,
	-1435599 when 7040,
	-1434398 when 7041,
	-1433196 when 7042,
	-1431993 when 7043,
	-1430790 when 7044,
	-1429585 when 7045,
	-1428379 when 7046,
	-1427173 when 7047,
	-1425966 when 7048,
	-1424757 when 7049,
	-1423548 when 7050,
	-1422338 when 7051,
	-1421128 when 7052,
	-1419916 when 7053,
	-1418703 when 7054,
	-1417490 when 7055,
	-1416276 when 7056,
	-1415060 when 7057,
	-1413844 when 7058,
	-1412627 when 7059,
	-1411410 when 7060,
	-1410191 when 7061,
	-1408971 when 7062,
	-1407751 when 7063,
	-1406530 when 7064,
	-1405307 when 7065,
	-1404084 when 7066,
	-1402861 when 7067,
	-1401636 when 7068,
	-1400410 when 7069,
	-1399184 when 7070,
	-1397956 when 7071,
	-1396728 when 7072,
	-1395499 when 7073,
	-1394269 when 7074,
	-1393038 when 7075,
	-1391807 when 7076,
	-1390574 when 7077,
	-1389341 when 7078,
	-1388107 when 7079,
	-1386872 when 7080,
	-1385636 when 7081,
	-1384399 when 7082,
	-1383161 when 7083,
	-1381923 when 7084,
	-1380683 when 7085,
	-1379443 when 7086,
	-1378202 when 7087,
	-1376960 when 7088,
	-1375717 when 7089,
	-1374474 when 7090,
	-1373229 when 7091,
	-1371984 when 7092,
	-1370738 when 7093,
	-1369491 when 7094,
	-1368243 when 7095,
	-1366994 when 7096,
	-1365745 when 7097,
	-1364495 when 7098,
	-1363243 when 7099,
	-1361991 when 7100,
	-1360738 when 7101,
	-1359485 when 7102,
	-1358230 when 7103,
	-1356975 when 7104,
	-1355718 when 7105,
	-1354461 when 7106,
	-1353203 when 7107,
	-1351945 when 7108,
	-1350685 when 7109,
	-1349425 when 7110,
	-1348164 when 7111,
	-1346901 when 7112,
	-1345639 when 7113,
	-1344375 when 7114,
	-1343110 when 7115,
	-1341845 when 7116,
	-1340579 when 7117,
	-1339312 when 7118,
	-1338044 when 7119,
	-1336775 when 7120,
	-1335505 when 7121,
	-1334235 when 7122,
	-1332964 when 7123,
	-1331692 when 7124,
	-1330419 when 7125,
	-1329146 when 7126,
	-1327871 when 7127,
	-1326596 when 7128,
	-1325320 when 7129,
	-1324043 when 7130,
	-1322765 when 7131,
	-1321487 when 7132,
	-1320207 when 7133,
	-1318927 when 7134,
	-1317646 when 7135,
	-1316364 when 7136,
	-1315082 when 7137,
	-1313798 when 7138,
	-1312514 when 7139,
	-1311229 when 7140,
	-1309943 when 7141,
	-1308656 when 7142,
	-1307369 when 7143,
	-1306081 when 7144,
	-1304792 when 7145,
	-1303502 when 7146,
	-1302211 when 7147,
	-1300920 when 7148,
	-1299627 when 7149,
	-1298334 when 7150,
	-1297040 when 7151,
	-1295746 when 7152,
	-1294450 when 7153,
	-1293154 when 7154,
	-1291857 when 7155,
	-1290559 when 7156,
	-1289260 when 7157,
	-1287961 when 7158,
	-1286660 when 7159,
	-1285359 when 7160,
	-1284057 when 7161,
	-1282755 when 7162,
	-1281451 when 7163,
	-1280147 when 7164,
	-1278842 when 7165,
	-1277536 when 7166,
	-1276230 when 7167,
	-1274922 when 7168,
	-1273614 when 7169,
	-1272305 when 7170,
	-1270995 when 7171,
	-1269685 when 7172,
	-1268374 when 7173,
	-1267061 when 7174,
	-1265749 when 7175,
	-1264435 when 7176,
	-1263120 when 7177,
	-1261805 when 7178,
	-1260489 when 7179,
	-1259172 when 7180,
	-1257855 when 7181,
	-1256537 when 7182,
	-1255218 when 7183,
	-1253898 when 7184,
	-1252577 when 7185,
	-1251256 when 7186,
	-1249933 when 7187,
	-1248610 when 7188,
	-1247287 when 7189,
	-1245962 when 7190,
	-1244637 when 7191,
	-1243311 when 7192,
	-1241984 when 7193,
	-1240656 when 7194,
	-1239328 when 7195,
	-1237999 when 7196,
	-1236669 when 7197,
	-1235339 when 7198,
	-1234007 when 7199,
	-1232675 when 7200,
	-1231342 when 7201,
	-1230008 when 7202,
	-1228674 when 7203,
	-1227339 when 7204,
	-1226003 when 7205,
	-1224666 when 7206,
	-1223329 when 7207,
	-1221991 when 7208,
	-1220652 when 7209,
	-1219312 when 7210,
	-1217971 when 7211,
	-1216630 when 7212,
	-1215288 when 7213,
	-1213945 when 7214,
	-1212602 when 7215,
	-1211258 when 7216,
	-1209913 when 7217,
	-1208567 when 7218,
	-1207221 when 7219,
	-1205873 when 7220,
	-1204525 when 7221,
	-1203177 when 7222,
	-1201827 when 7223,
	-1200477 when 7224,
	-1199126 when 7225,
	-1197775 when 7226,
	-1196422 when 7227,
	-1195069 when 7228,
	-1193715 when 7229,
	-1192361 when 7230,
	-1191005 when 7231,
	-1189649 when 7232,
	-1188292 when 7233,
	-1186935 when 7234,
	-1185577 when 7235,
	-1184218 when 7236,
	-1182858 when 7237,
	-1181497 when 7238,
	-1180136 when 7239,
	-1178774 when 7240,
	-1177412 when 7241,
	-1176048 when 7242,
	-1174684 when 7243,
	-1173319 when 7244,
	-1171954 when 7245,
	-1170588 when 7246,
	-1169221 when 7247,
	-1167853 when 7248,
	-1166484 when 7249,
	-1165115 when 7250,
	-1163745 when 7251,
	-1162375 when 7252,
	-1161003 when 7253,
	-1159631 when 7254,
	-1158259 when 7255,
	-1156885 when 7256,
	-1155511 when 7257,
	-1154136 when 7258,
	-1152761 when 7259,
	-1151384 when 7260,
	-1150007 when 7261,
	-1148630 when 7262,
	-1147251 when 7263,
	-1145872 when 7264,
	-1144492 when 7265,
	-1143112 when 7266,
	-1141730 when 7267,
	-1140348 when 7268,
	-1138966 when 7269,
	-1137582 when 7270,
	-1136198 when 7271,
	-1134814 when 7272,
	-1133428 when 7273,
	-1132042 when 7274,
	-1130655 when 7275,
	-1129267 when 7276,
	-1127879 when 7277,
	-1126490 when 7278,
	-1125101 when 7279,
	-1123710 when 7280,
	-1122319 when 7281,
	-1120927 when 7282,
	-1119535 when 7283,
	-1118142 when 7284,
	-1116748 when 7285,
	-1115354 when 7286,
	-1113958 when 7287,
	-1112563 when 7288,
	-1111166 when 7289,
	-1109769 when 7290,
	-1108371 when 7291,
	-1106972 when 7292,
	-1105573 when 7293,
	-1104173 when 7294,
	-1102772 when 7295,
	-1101371 when 7296,
	-1099969 when 7297,
	-1098566 when 7298,
	-1097163 when 7299,
	-1095759 when 7300,
	-1094354 when 7301,
	-1092949 when 7302,
	-1091543 when 7303,
	-1090136 when 7304,
	-1088729 when 7305,
	-1087320 when 7306,
	-1085912 when 7307,
	-1084502 when 7308,
	-1083092 when 7309,
	-1081681 when 7310,
	-1080270 when 7311,
	-1078858 when 7312,
	-1077445 when 7313,
	-1076032 when 7314,
	-1074618 when 7315,
	-1073203 when 7316,
	-1071787 when 7317,
	-1070371 when 7318,
	-1068955 when 7319,
	-1067537 when 7320,
	-1066119 when 7321,
	-1064700 when 7322,
	-1063281 when 7323,
	-1061861 when 7324,
	-1060440 when 7325,
	-1059019 when 7326,
	-1057597 when 7327,
	-1056174 when 7328,
	-1054751 when 7329,
	-1053327 when 7330,
	-1051903 when 7331,
	-1050477 when 7332,
	-1049051 when 7333,
	-1047625 when 7334,
	-1046198 when 7335,
	-1044770 when 7336,
	-1043341 when 7337,
	-1041912 when 7338,
	-1040483 when 7339,
	-1039052 when 7340,
	-1037621 when 7341,
	-1036189 when 7342,
	-1034757 when 7343,
	-1033324 when 7344,
	-1031891 when 7345,
	-1030456 when 7346,
	-1029021 when 7347,
	-1027586 when 7348,
	-1026150 when 7349,
	-1024713 when 7350,
	-1023276 when 7351,
	-1021838 when 7352,
	-1020399 when 7353,
	-1018960 when 7354,
	-1017520 when 7355,
	-1016079 when 7356,
	-1014638 when 7357,
	-1013196 when 7358,
	-1011754 when 7359,
	-1010311 when 7360,
	-1008867 when 7361,
	-1007423 when 7362,
	-1005978 when 7363,
	-1004532 when 7364,
	-1003086 when 7365,
	-1001639 when 7366,
	-1000192 when 7367,
	-998744 when 7368,
	-997295 when 7369,
	-995846 when 7370,
	-994396 when 7371,
	-992946 when 7372,
	-991495 when 7373,
	-990043 when 7374,
	-988591 when 7375,
	-987138 when 7376,
	-985684 when 7377,
	-984230 when 7378,
	-982775 when 7379,
	-981320 when 7380,
	-979864 when 7381,
	-978407 when 7382,
	-976950 when 7383,
	-975493 when 7384,
	-974034 when 7385,
	-972575 when 7386,
	-971116 when 7387,
	-969655 when 7388,
	-968195 when 7389,
	-966733 when 7390,
	-965271 when 7391,
	-963809 when 7392,
	-962346 when 7393,
	-960882 when 7394,
	-959418 when 7395,
	-957953 when 7396,
	-956487 when 7397,
	-955021 when 7398,
	-953554 when 7399,
	-952087 when 7400,
	-950619 when 7401,
	-949151 when 7402,
	-947682 when 7403,
	-946212 when 7404,
	-944742 when 7405,
	-943271 when 7406,
	-941800 when 7407,
	-940328 when 7408,
	-938855 when 7409,
	-937382 when 7410,
	-935908 when 7411,
	-934434 when 7412,
	-932959 when 7413,
	-931484 when 7414,
	-930008 when 7415,
	-928531 when 7416,
	-927054 when 7417,
	-925576 when 7418,
	-924098 when 7419,
	-922619 when 7420,
	-921140 when 7421,
	-919660 when 7422,
	-918179 when 7423,
	-916698 when 7424,
	-915217 when 7425,
	-913734 when 7426,
	-912251 when 7427,
	-910768 when 7428,
	-909284 when 7429,
	-907800 when 7430,
	-906315 when 7431,
	-904829 when 7432,
	-903343 when 7433,
	-901856 when 7434,
	-900369 when 7435,
	-898881 when 7436,
	-897392 when 7437,
	-895903 when 7438,
	-894414 when 7439,
	-892924 when 7440,
	-891433 when 7441,
	-889942 when 7442,
	-888450 when 7443,
	-886958 when 7444,
	-885465 when 7445,
	-883972 when 7446,
	-882478 when 7447,
	-880984 when 7448,
	-879489 when 7449,
	-877993 when 7450,
	-876497 when 7451,
	-875000 when 7452,
	-873503 when 7453,
	-872006 when 7454,
	-870507 when 7455,
	-869009 when 7456,
	-867509 when 7457,
	-866009 when 7458,
	-864509 when 7459,
	-863008 when 7460,
	-861507 when 7461,
	-860005 when 7462,
	-858502 when 7463,
	-856999 when 7464,
	-855496 when 7465,
	-853992 when 7466,
	-852487 when 7467,
	-850982 when 7468,
	-849476 when 7469,
	-847970 when 7470,
	-846463 when 7471,
	-844956 when 7472,
	-843448 when 7473,
	-841940 when 7474,
	-840431 when 7475,
	-838922 when 7476,
	-837412 when 7477,
	-835902 when 7478,
	-834391 when 7479,
	-832879 when 7480,
	-831368 when 7481,
	-829855 when 7482,
	-828342 when 7483,
	-826829 when 7484,
	-825315 when 7485,
	-823800 when 7486,
	-822286 when 7487,
	-820770 when 7488,
	-819254 when 7489,
	-817738 when 7490,
	-816221 when 7491,
	-814703 when 7492,
	-813185 when 7493,
	-811667 when 7494,
	-810148 when 7495,
	-808628 when 7496,
	-807108 when 7497,
	-805588 when 7498,
	-804067 when 7499,
	-802545 when 7500,
	-801023 when 7501,
	-799501 when 7502,
	-797978 when 7503,
	-796454 when 7504,
	-794931 when 7505,
	-793406 when 7506,
	-791881 when 7507,
	-790356 when 7508,
	-788830 when 7509,
	-787304 when 7510,
	-785777 when 7511,
	-784249 when 7512,
	-782721 when 7513,
	-781193 when 7514,
	-779664 when 7515,
	-778135 when 7516,
	-776605 when 7517,
	-775075 when 7518,
	-773544 when 7519,
	-772013 when 7520,
	-770481 when 7521,
	-768949 when 7522,
	-767417 when 7523,
	-765884 when 7524,
	-764350 when 7525,
	-762816 when 7526,
	-761281 when 7527,
	-759747 when 7528,
	-758211 when 7529,
	-756675 when 7530,
	-755139 when 7531,
	-753602 when 7532,
	-752065 when 7533,
	-750527 when 7534,
	-748989 when 7535,
	-747450 when 7536,
	-745911 when 7537,
	-744371 when 7538,
	-742831 when 7539,
	-741290 when 7540,
	-739749 when 7541,
	-738208 when 7542,
	-736666 when 7543,
	-735124 when 7544,
	-733581 when 7545,
	-732038 when 7546,
	-730494 when 7547,
	-728950 when 7548,
	-727405 when 7549,
	-725860 when 7550,
	-724315 when 7551,
	-722769 when 7552,
	-721222 when 7553,
	-719675 when 7554,
	-718128 when 7555,
	-716580 when 7556,
	-715032 when 7557,
	-713483 when 7558,
	-711934 when 7559,
	-710385 when 7560,
	-708835 when 7561,
	-707285 when 7562,
	-705734 when 7563,
	-704183 when 7564,
	-702631 when 7565,
	-701079 when 7566,
	-699526 when 7567,
	-697973 when 7568,
	-696420 when 7569,
	-694866 when 7570,
	-693312 when 7571,
	-691757 when 7572,
	-690202 when 7573,
	-688646 when 7574,
	-687090 when 7575,
	-685534 when 7576,
	-683977 when 7577,
	-682420 when 7578,
	-680862 when 7579,
	-679304 when 7580,
	-677746 when 7581,
	-676187 when 7582,
	-674627 when 7583,
	-673068 when 7584,
	-671507 when 7585,
	-669947 when 7586,
	-668386 when 7587,
	-666824 when 7588,
	-665263 when 7589,
	-663700 when 7590,
	-662138 when 7591,
	-660575 when 7592,
	-659011 when 7593,
	-657447 when 7594,
	-655883 when 7595,
	-654318 when 7596,
	-652753 when 7597,
	-651188 when 7598,
	-649622 when 7599,
	-648056 when 7600,
	-646489 when 7601,
	-644922 when 7602,
	-643354 when 7603,
	-641786 when 7604,
	-640218 when 7605,
	-638650 when 7606,
	-637080 when 7607,
	-635511 when 7608,
	-633941 when 7609,
	-632371 when 7610,
	-630800 when 7611,
	-629229 when 7612,
	-627658 when 7613,
	-626086 when 7614,
	-624514 when 7615,
	-622941 when 7616,
	-621368 when 7617,
	-619795 when 7618,
	-618221 when 7619,
	-616647 when 7620,
	-615073 when 7621,
	-613498 when 7622,
	-611923 when 7623,
	-610347 when 7624,
	-608771 when 7625,
	-607195 when 7626,
	-605618 when 7627,
	-604041 when 7628,
	-602463 when 7629,
	-600886 when 7630,
	-599307 when 7631,
	-597729 when 7632,
	-596150 when 7633,
	-594570 when 7634,
	-592991 when 7635,
	-591411 when 7636,
	-589830 when 7637,
	-588249 when 7638,
	-586668 when 7639,
	-585087 when 7640,
	-583505 when 7641,
	-581923 when 7642,
	-580340 when 7643,
	-578757 when 7644,
	-577174 when 7645,
	-575590 when 7646,
	-574006 when 7647,
	-572422 when 7648,
	-570837 when 7649,
	-569252 when 7650,
	-567666 when 7651,
	-566081 when 7652,
	-564495 when 7653,
	-562908 when 7654,
	-561321 when 7655,
	-559734 when 7656,
	-558147 when 7657,
	-556559 when 7658,
	-554970 when 7659,
	-553382 when 7660,
	-551793 when 7661,
	-550204 when 7662,
	-548614 when 7663,
	-547024 when 7664,
	-545434 when 7665,
	-543843 when 7666,
	-542253 when 7667,
	-540661 when 7668,
	-539070 when 7669,
	-537478 when 7670,
	-535886 when 7671,
	-534293 when 7672,
	-532700 when 7673,
	-531107 when 7674,
	-529513 when 7675,
	-527919 when 7676,
	-526325 when 7677,
	-524731 when 7678,
	-523136 when 7679,
	-521540 when 7680,
	-519945 when 7681,
	-518349 when 7682,
	-516753 when 7683,
	-515157 when 7684,
	-513560 when 7685,
	-511963 when 7686,
	-510365 when 7687,
	-508767 when 7688,
	-507169 when 7689,
	-505571 when 7690,
	-503972 when 7691,
	-502373 when 7692,
	-500774 when 7693,
	-499174 when 7694,
	-497575 when 7695,
	-495974 when 7696,
	-494374 when 7697,
	-492773 when 7698,
	-491172 when 7699,
	-489570 when 7700,
	-487969 when 7701,
	-486367 when 7702,
	-484764 when 7703,
	-483162 when 7704,
	-481559 when 7705,
	-479955 when 7706,
	-478352 when 7707,
	-476748 when 7708,
	-475144 when 7709,
	-473540 when 7710,
	-471935 when 7711,
	-470330 when 7712,
	-468725 when 7713,
	-467119 when 7714,
	-465513 when 7715,
	-463907 when 7716,
	-462301 when 7717,
	-460694 when 7718,
	-459087 when 7719,
	-457480 when 7720,
	-455872 when 7721,
	-454264 when 7722,
	-452656 when 7723,
	-451048 when 7724,
	-449439 when 7725,
	-447830 when 7726,
	-446221 when 7727,
	-444611 when 7728,
	-443001 when 7729,
	-441391 when 7730,
	-439781 when 7731,
	-438170 when 7732,
	-436559 when 7733,
	-434948 when 7734,
	-433337 when 7735,
	-431725 when 7736,
	-430113 when 7737,
	-428501 when 7738,
	-426889 when 7739,
	-425276 when 7740,
	-423663 when 7741,
	-422050 when 7742,
	-420436 when 7743,
	-418822 when 7744,
	-417208 when 7745,
	-415594 when 7746,
	-413979 when 7747,
	-412364 when 7748,
	-410749 when 7749,
	-409134 when 7750,
	-407518 when 7751,
	-405903 when 7752,
	-404287 when 7753,
	-402670 when 7754,
	-401054 when 7755,
	-399437 when 7756,
	-397820 when 7757,
	-396202 when 7758,
	-394585 when 7759,
	-392967 when 7760,
	-391349 when 7761,
	-389731 when 7762,
	-388112 when 7763,
	-386493 when 7764,
	-384874 when 7765,
	-383255 when 7766,
	-381636 when 7767,
	-380016 when 7768,
	-378396 when 7769,
	-376776 when 7770,
	-375155 when 7771,
	-373535 when 7772,
	-371914 when 7773,
	-370293 when 7774,
	-368672 when 7775,
	-367050 when 7776,
	-365428 when 7777,
	-363806 when 7778,
	-362184 when 7779,
	-360561 when 7780,
	-358939 when 7781,
	-357316 when 7782,
	-355693 when 7783,
	-354069 when 7784,
	-352446 when 7785,
	-350822 when 7786,
	-349198 when 7787,
	-347574 when 7788,
	-345949 when 7789,
	-344325 when 7790,
	-342700 when 7791,
	-341075 when 7792,
	-339450 when 7793,
	-337824 when 7794,
	-336198 when 7795,
	-334573 when 7796,
	-332946 when 7797,
	-331320 when 7798,
	-329694 when 7799,
	-328067 when 7800,
	-326440 when 7801,
	-324813 when 7802,
	-323185 when 7803,
	-321558 when 7804,
	-319930 when 7805,
	-318302 when 7806,
	-316674 when 7807,
	-315046 when 7808,
	-313417 when 7809,
	-311789 when 7810,
	-310160 when 7811,
	-308531 when 7812,
	-306901 when 7813,
	-305272 when 7814,
	-303642 when 7815,
	-302013 when 7816,
	-300382 when 7817,
	-298752 when 7818,
	-297122 when 7819,
	-295491 when 7820,
	-293861 when 7821,
	-292230 when 7822,
	-290598 when 7823,
	-288967 when 7824,
	-287336 when 7825,
	-285704 when 7826,
	-284072 when 7827,
	-282440 when 7828,
	-280808 when 7829,
	-279176 when 7830,
	-277543 when 7831,
	-275910 when 7832,
	-274278 when 7833,
	-272645 when 7834,
	-271011 when 7835,
	-269378 when 7836,
	-267744 when 7837,
	-266111 when 7838,
	-264477 when 7839,
	-262843 when 7840,
	-261209 when 7841,
	-259574 when 7842,
	-257940 when 7843,
	-256305 when 7844,
	-254670 when 7845,
	-253035 when 7846,
	-251400 when 7847,
	-249765 when 7848,
	-248129 when 7849,
	-246494 when 7850,
	-244858 when 7851,
	-243222 when 7852,
	-241586 when 7853,
	-239950 when 7854,
	-238313 when 7855,
	-236677 when 7856,
	-235040 when 7857,
	-233404 when 7858,
	-231767 when 7859,
	-230130 when 7860,
	-228492 when 7861,
	-226855 when 7862,
	-225217 when 7863,
	-223580 when 7864,
	-221942 when 7865,
	-220304 when 7866,
	-218666 when 7867,
	-217028 when 7868,
	-215390 when 7869,
	-213751 when 7870,
	-212112 when 7871,
	-210474 when 7872,
	-208835 when 7873,
	-207196 when 7874,
	-205557 when 7875,
	-203918 when 7876,
	-202278 when 7877,
	-200639 when 7878,
	-198999 when 7879,
	-197359 when 7880,
	-195720 when 7881,
	-194080 when 7882,
	-192440 when 7883,
	-190799 when 7884,
	-189159 when 7885,
	-187519 when 7886,
	-185878 when 7887,
	-184237 when 7888,
	-182597 when 7889,
	-180956 when 7890,
	-179315 when 7891,
	-177673 when 7892,
	-176032 when 7893,
	-174391 when 7894,
	-172749 when 7895,
	-171108 when 7896,
	-169466 when 7897,
	-167824 when 7898,
	-166183 when 7899,
	-164541 when 7900,
	-162899 when 7901,
	-161256 when 7902,
	-159614 when 7903,
	-157972 when 7904,
	-156329 when 7905,
	-154687 when 7906,
	-153044 when 7907,
	-151401 when 7908,
	-149758 when 7909,
	-148116 when 7910,
	-146472 when 7911,
	-144829 when 7912,
	-143186 when 7913,
	-141543 when 7914,
	-139899 when 7915,
	-138256 when 7916,
	-136612 when 7917,
	-134969 when 7918,
	-133325 when 7919,
	-131681 when 7920,
	-130037 when 7921,
	-128393 when 7922,
	-126749 when 7923,
	-125105 when 7924,
	-123461 when 7925,
	-121817 when 7926,
	-120172 when 7927,
	-118528 when 7928,
	-116883 when 7929,
	-115239 when 7930,
	-113594 when 7931,
	-111950 when 7932,
	-110305 when 7933,
	-108660 when 7934,
	-107015 when 7935,
	-105370 when 7936,
	-103725 when 7937,
	-102080 when 7938,
	-100435 when 7939,
	-98789 when 7940,
	-97144 when 7941,
	-95499 when 7942,
	-93853 when 7943,
	-92208 when 7944,
	-90562 when 7945,
	-88917 when 7946,
	-87271 when 7947,
	-85625 when 7948,
	-83980 when 7949,
	-82334 when 7950,
	-80688 when 7951,
	-79042 when 7952,
	-77396 when 7953,
	-75750 when 7954,
	-74104 when 7955,
	-72458 when 7956,
	-70812 when 7957,
	-69166 when 7958,
	-67519 when 7959,
	-65873 when 7960,
	-64227 when 7961,
	-62580 when 7962,
	-60934 when 7963,
	-59288 when 7964,
	-57641 when 7965,
	-55995 when 7966,
	-54348 when 7967,
	-52702 when 7968,
	-51055 when 7969,
	-49408 when 7970,
	-47762 when 7971,
	-46115 when 7972,
	-44468 when 7973,
	-42822 when 7974,
	-41175 when 7975,
	-39528 when 7976,
	-37881 when 7977,
	-36234 when 7978,
	-34588 when 7979,
	-32941 when 7980,
	-31294 when 7981,
	-29647 when 7982,
	-28000 when 7983,
	-26353 when 7984,
	-24706 when 7985,
	-23059 when 7986,
	-21412 when 7987,
	-19765 when 7988,
	-18118 when 7989,
	-16471 when 7990,
	-14824 when 7991,
	-13177 when 7992,
	-11530 when 7993,
	-9883 when 7994,
	-8235 when 7995,
	-6588 when 7996,
	-4941 when 7997,
	-3294 when 7998,
	-1647 when 7999,					
							0 when others;

end rtl;