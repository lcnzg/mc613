library ieee;
use ieee.std_logic_1164.all;

entity sine_wave is
	port (
		indice: in integer range 0 to 4095;
		amplitude: out integer range -2097152 to 2097152
);
end sine_wave;

architecture rtl of sine_wave is

begin

	with indice select
		amplitude <=
			0 when 0,
			3217 when 1,
			6434 when 2,
			9651 when 3,
			12868 when 4,
			16085 when 5,
			19302 when 6,
			22519 when 7,
			25735 when 8,
			28952 when 9,
			32169 when 10,
			35385 when 11,
			38602 when 12,
			41818 when 13,
			45034 when 14,
			48251 when 15,
			51467 when 16,
			54683 when 17,
			57898 when 18,
			61114 when 19,
			64330 when 20,
			67545 when 21,
			70760 when 22,
			73975 when 23,
			77190 when 24,
			80405 when 25,
			83620 when 26,
			86834 when 27,
			90048 when 28,
			93262 when 29,
			96476 when 30,
			99689 when 31,
			102902 when 32,
			106115 when 33,
			109328 when 34,
			112541 when 35,
			115753 when 36,
			118965 when 37,
			122176 when 38,
			125388 when 39,
			128599 when 40,
			131810 when 41,
			135020 when 42,
			138230 when 43,
			141440 when 44,
			144650 when 45,
			147859 when 46,
			151068 when 47,
			154276 when 48,
			157484 when 49,
			160692 when 50,
			163899 when 51,
			167106 when 52,
			170313 when 53,
			173519 when 54,
			176725 when 55,
			179930 when 56,
			183135 when 57,
			186339 when 58,
			189543 when 59,
			192747 when 60,
			195950 when 61,
			199153 when 62,
			202355 when 63,
			205557 when 64,
			208758 when 65,
			211959 when 66,
			215159 when 67,
			218359 when 68,
			221558 when 69,
			224757 when 70,
			227955 when 71,
			231153 when 72,
			234350 when 73,
			237546 when 74,
			240742 when 75,
			243938 when 76,
			247133 when 77,
			250327 when 78,
			253521 when 79,
			256714 when 80,
			259906 when 81,
			263098 when 82,
			266289 when 83,
			269480 when 84,
			272670 when 85,
			275859 when 86,
			279048 when 87,
			282236 when 88,
			285424 when 89,
			288610 when 90,
			291796 when 91,
			294982 when 92,
			298166 when 93,
			301350 when 94,
			304534 when 95,
			307716 when 96,
			310898 when 97,
			314079 when 98,
			317259 when 99,
			320439 when 100,
			323618 when 101,
			326796 when 102,
			329973 when 103,
			333150 when 104,
			336325 when 105,
			339500 when 106,
			342675 when 107,
			345848 when 108,
			349020 when 109,
			352192 when 110,
			355363 when 111,
			358533 when 112,
			361702 when 113,
			364871 when 114,
			368038 when 115,
			371205 when 116,
			374371 when 117,
			377535 when 118,
			380699 when 119,
			383862 when 120,
			387025 when 121,
			390186 when 122,
			393346 when 123,
			396506 when 124,
			399664 when 125,
			402822 when 126,
			405978 when 127,
			409134 when 128,
			412289 when 129,
			415442 when 130,
			418595 when 131,
			421747 when 132,
			424898 when 133,
			428048 when 134,
			431196 when 135,
			434344 when 136,
			437491 when 137,
			440636 when 138,
			443781 when 139,
			446925 when 140,
			450067 when 141,
			453209 when 142,
			456349 when 143,
			459489 when 144,
			462627 when 145,
			465764 when 146,
			468900 when 147,
			472035 when 148,
			475169 when 149,
			478302 when 150,
			481433 when 151,
			484564 when 152,
			487693 when 153,
			490822 when 154,
			493949 when 155,
			497075 when 156,
			500199 when 157,
			503323 when 158,
			506445 when 159,
			509566 when 160,
			512686 when 161,
			515805 when 162,
			518923 when 163,
			522039 when 164,
			525154 when 165,
			528268 when 166,
			531381 when 167,
			534492 when 168,
			537602 when 169,
			540711 when 170,
			543819 when 171,
			546925 when 172,
			550030 when 173,
			553134 when 174,
			556236 when 175,
			559337 when 176,
			562437 when 177,
			565535 when 178,
			568633 when 179,
			571728 when 180,
			574823 when 181,
			577916 when 182,
			581008 when 183,
			584098 when 184,
			587187 when 185,
			590275 when 186,
			593361 when 187,
			596446 when 188,
			599529 when 189,
			602611 when 190,
			605692 when 191,
			608771 when 192,
			611849 when 193,
			614925 when 194,
			618000 when 195,
			621073 when 196,
			624145 when 197,
			627216 when 198,
			630285 when 199,
			633352 when 200,
			636418 when 201,
			639483 when 202,
			642546 when 203,
			645607 when 204,
			648667 when 205,
			651726 when 206,
			654783 when 207,
			657838 when 208,
			660892 when 209,
			663944 when 210,
			666995 when 211,
			670044 when 212,
			673092 when 213,
			676138 when 214,
			679182 when 215,
			682225 when 216,
			685266 when 217,
			688306 when 218,
			691344 when 219,
			694380 when 220,
			697415 when 221,
			700448 when 222,
			703479 when 223,
			706509 when 224,
			709537 when 225,
			712564 when 226,
			715589 when 227,
			718612 when 228,
			721633 when 229,
			724653 when 230,
			727671 when 231,
			730687 when 232,
			733701 when 233,
			736714 when 234,
			739725 when 235,
			742735 when 236,
			745742 when 237,
			748748 when 238,
			751752 when 239,
			754755 when 240,
			757755 when 241,
			760754 when 242,
			763751 when 243,
			766746 when 244,
			769739 when 245,
			772731 when 246,
			775721 when 247,
			778709 when 248,
			781695 when 249,
			784679 when 250,
			787661 when 251,
			790642 when 252,
			793621 when 253,
			796597 when 254,
			799572 when 255,
			802545 when 256,
			805516 when 257,
			808486 when 258,
			811453 when 259,
			814419 when 260,
			817382 when 261,
			820344 when 262,
			823303 when 263,
			826261 when 264,
			829217 when 265,
			832171 when 266,
			835123 when 267,
			838073 when 268,
			841021 when 269,
			843967 when 270,
			846911 when 271,
			849853 when 272,
			852793 when 273,
			855731 when 274,
			858667 when 275,
			861601 when 276,
			864533 when 277,
			867462 when 278,
			870390 when 279,
			873316 when 280,
			876240 when 281,
			879162 when 282,
			882081 when 283,
			884999 when 284,
			887914 when 285,
			890828 when 286,
			893739 when 287,
			896648 when 288,
			899555 when 289,
			902460 when 290,
			905363 when 291,
			908264 when 292,
			911162 when 293,
			914059 when 294,
			916953 when 295,
			919845 when 296,
			922735 when 297,
			925623 when 298,
			928508 when 299,
			931392 when 300,
			934273 when 301,
			937152 when 302,
			940029 when 303,
			942903 when 304,
			945776 when 305,
			948646 when 306,
			951514 when 307,
			954379 when 308,
			957243 when 309,
			960104 when 310,
			962963 when 311,
			965820 when 312,
			968674 when 313,
			971526 when 314,
			974376 when 315,
			977224 when 316,
			980069 when 317,
			982912 when 318,
			985752 when 319,
			988591 when 320,
			991427 when 321,
			994260 when 322,
			997092 when 323,
			999920 when 324,
			1002747 when 325,
			1005571 when 326,
			1008393 when 327,
			1011213 when 328,
			1014030 when 329,
			1016845 when 330,
			1019657 when 331,
			1022467 when 332,
			1025274 when 333,
			1028079 when 334,
			1030882 when 335,
			1033682 when 336,
			1036480 when 337,
			1039276 when 338,
			1042069 when 339,
			1044859 when 340,
			1047647 when 341,
			1050433 when 342,
			1053216 when 343,
			1055997 when 344,
			1058775 when 345,
			1061550 when 346,
			1064323 when 347,
			1067094 when 348,
			1069862 when 349,
			1072628 when 350,
			1075391 when 351,
			1078152 when 352,
			1080910 when 353,
			1083665 when 354,
			1086418 when 355,
			1089168 when 356,
			1091916 when 357,
			1094662 when 358,
			1097404 when 359,
			1100144 when 360,
			1102882 when 361,
			1105617 when 362,
			1108349 when 363,
			1111079 when 364,
			1113806 when 365,
			1116530 when 366,
			1119252 when 367,
			1121971 when 368,
			1124688 when 369,
			1127402 when 370,
			1130113 when 371,
			1132822 when 372,
			1135528 when 373,
			1138231 when 374,
			1140931 when 375,
			1143629 when 376,
			1146325 when 377,
			1149017 when 378,
			1151707 when 379,
			1154394 when 380,
			1157078 when 381,
			1159760 when 382,
			1162439 when 383,
			1165115 when 384,
			1167789 when 385,
			1170459 when 386,
			1173127 when 387,
			1175793 when 388,
			1178455 when 389,
			1181115 when 390,
			1183772 when 391,
			1186426 when 392,
			1189077 when 393,
			1191725 when 394,
			1194371 when 395,
			1197014 when 396,
			1199654 when 397,
			1202291 when 398,
			1204926 when 399,
			1207557 when 400,
			1210186 when 401,
			1212812 when 402,
			1215435 when 403,
			1218055 when 404,
			1220672 when 405,
			1223287 when 406,
			1225898 when 407,
			1228507 when 408,
			1231113 when 409,
			1233716 when 410,
			1236316 when 411,
			1238913 when 412,
			1241507 when 413,
			1244098 when 414,
			1246687 when 415,
			1249272 when 416,
			1251854 when 417,
			1254434 when 418,
			1257010 when 419,
			1259584 when 420,
			1262155 when 421,
			1264722 when 422,
			1267287 when 423,
			1269849 when 424,
			1272407 when 425,
			1274963 when 426,
			1277516 when 427,
			1280066 when 428,
			1282612 when 429,
			1285156 when 430,
			1287697 when 431,
			1290234 when 432,
			1292769 when 433,
			1295300 when 434,
			1297829 when 435,
			1300354 when 436,
			1302877 when 437,
			1305396 when 438,
			1307912 when 439,
			1310425 when 440,
			1312935 when 441,
			1315442 when 442,
			1317946 when 443,
			1320447 when 444,
			1322945 when 445,
			1325439 when 446,
			1327931 when 447,
			1330419 when 448,
			1332904 when 449,
			1335386 when 450,
			1337865 when 451,
			1340341 when 452,
			1342814 when 453,
			1345283 when 454,
			1347749 when 455,
			1350213 when 456,
			1352673 when 457,
			1355129 when 458,
			1357583 when 459,
			1360033 when 460,
			1362480 when 461,
			1364924 when 462,
			1367365 when 463,
			1369803 when 464,
			1372237 when 465,
			1374668 when 466,
			1377096 when 467,
			1379521 when 468,
			1381942 when 469,
			1384360 when 470,
			1386775 when 471,
			1389187 when 472,
			1391595 when 473,
			1394000 when 474,
			1396402 when 475,
			1398800 when 476,
			1401195 when 477,
			1403587 when 478,
			1405976 when 479,
			1408361 when 480,
			1410743 when 481,
			1413122 when 482,
			1415497 when 483,
			1417869 when 484,
			1420238 when 485,
			1422603 when 486,
			1424965 when 487,
			1427324 when 488,
			1429679 when 489,
			1432031 when 490,
			1434379 when 491,
			1436725 when 492,
			1439066 when 493,
			1441405 when 494,
			1443740 when 495,
			1446071 when 496,
			1448400 when 497,
			1450724 when 498,
			1453046 when 499,
			1455364 when 500,
			1457678 when 501,
			1459989 when 502,
			1462297 when 503,
			1464601 when 504,
			1466902 when 505,
			1469199 when 506,
			1471493 when 507,
			1473784 when 508,
			1476070 when 509,
			1478354 when 510,
			1480634 when 511,
			1482910 when 512,
			1485183 when 513,
			1487453 when 514,
			1489719 when 515,
			1491981 when 516,
			1494240 when 517,
			1496496 when 518,
			1498748 when 519,
			1500996 when 520,
			1503241 when 521,
			1505483 when 522,
			1507720 when 523,
			1509955 when 524,
			1512185 when 525,
			1514413 when 526,
			1516636 when 527,
			1518856 when 528,
			1521073 when 529,
			1523286 when 530,
			1525495 when 531,
			1527701 when 532,
			1529903 when 533,
			1532101 when 534,
			1534296 when 535,
			1536487 when 536,
			1538675 when 537,
			1540859 when 538,
			1543040 when 539,
			1545216 when 540,
			1547390 when 541,
			1549559 when 542,
			1551725 when 543,
			1553887 when 544,
			1556046 when 545,
			1558201 when 546,
			1560352 when 547,
			1562499 when 548,
			1564643 when 549,
			1566784 when 550,
			1568920 when 551,
			1571053 when 552,
			1573182 when 553,
			1575307 when 554,
			1577429 when 555,
			1579547 when 556,
			1581662 when 557,
			1583772 when 558,
			1585879 when 559,
			1587982 when 560,
			1590081 when 561,
			1592177 when 562,
			1594269 when 563,
			1596357 when 564,
			1598441 when 565,
			1600522 when 566,
			1602599 when 567,
			1604672 when 568,
			1606741 when 569,
			1608807 when 570,
			1610869 when 571,
			1612927 when 572,
			1614981 when 573,
			1617031 when 574,
			1619078 when 575,
			1621120 when 576,
			1623159 when 577,
			1625194 when 578,
			1627226 when 579,
			1629253 when 580,
			1631277 when 581,
			1633297 when 582,
			1635313 when 583,
			1637325 when 584,
			1639333 when 585,
			1641337 when 586,
			1643338 when 587,
			1645334 when 588,
			1647327 when 589,
			1649316 when 590,
			1651301 when 591,
			1653282 when 592,
			1655260 when 593,
			1657233 when 594,
			1659202 when 595,
			1661168 when 596,
			1663130 when 597,
			1665087 when 598,
			1667041 when 599,
			1668991 when 600,
			1670937 when 601,
			1672879 when 602,
			1674817 when 603,
			1676751 when 604,
			1678681 when 605,
			1680608 when 606,
			1682530 when 607,
			1684448 when 608,
			1686363 when 609,
			1688273 when 610,
			1690180 when 611,
			1692082 when 612,
			1693980 when 613,
			1695875 when 614,
			1697765 when 615,
			1699652 when 616,
			1701534 when 617,
			1703413 when 618,
			1705287 when 619,
			1707158 when 620,
			1709024 when 621,
			1710887 when 622,
			1712745 when 623,
			1714600 when 624,
			1716450 when 625,
			1718296 when 626,
			1720139 when 627,
			1721977 when 628,
			1723811 when 629,
			1725641 when 630,
			1727467 when 631,
			1729289 when 632,
			1731107 when 633,
			1732921 when 634,
			1734731 when 635,
			1736536 when 636,
			1738338 when 637,
			1740135 when 638,
			1741929 when 639,
			1743718 when 640,
			1745503 when 641,
			1747284 when 642,
			1749061 when 643,
			1750834 when 644,
			1752603 when 645,
			1754368 when 646,
			1756128 when 647,
			1757885 when 648,
			1759637 when 649,
			1761385 when 650,
			1763129 when 651,
			1764869 when 652,
			1766604 when 653,
			1768336 when 654,
			1770063 when 655,
			1771786 when 656,
			1773505 when 657,
			1775220 when 658,
			1776931 when 659,
			1778637 when 660,
			1780340 when 661,
			1782038 when 662,
			1783732 when 663,
			1785421 when 664,
			1787107 when 665,
			1788788 when 666,
			1790465 when 667,
			1792138 when 668,
			1793807 when 669,
			1795471 when 670,
			1797131 when 671,
			1798787 when 672,
			1800439 when 673,
			1802087 when 674,
			1803730 when 675,
			1805369 when 676,
			1807004 when 677,
			1808634 when 678,
			1810260 when 679,
			1811882 when 680,
			1813500 when 681,
			1815114 when 682,
			1816723 when 683,
			1818328 when 684,
			1819928 when 685,
			1821525 when 686,
			1823117 when 687,
			1824705 when 688,
			1826288 when 689,
			1827867 when 690,
			1829442 when 691,
			1831013 when 692,
			1832579 when 693,
			1834141 when 694,
			1835699 when 695,
			1837252 when 696,
			1838801 when 697,
			1840346 when 698,
			1841886 when 699,
			1843422 when 700,
			1844954 when 701,
			1846481 when 702,
			1848004 when 703,
			1849523 when 704,
			1851037 when 705,
			1852547 when 706,
			1854053 when 707,
			1855554 when 708,
			1857051 when 709,
			1858543 when 710,
			1860031 when 711,
			1861515 when 712,
			1862995 when 713,
			1864470 when 714,
			1865940 when 715,
			1867406 when 716,
			1868868 when 717,
			1870326 when 718,
			1871779 when 719,
			1873227 when 720,
			1874671 when 721,
			1876111 when 722,
			1877546 when 723,
			1878977 when 724,
			1880404 when 725,
			1881826 when 726,
			1883244 when 727,
			1884657 when 728,
			1886066 when 729,
			1887470 when 730,
			1888870 when 731,
			1890266 when 732,
			1891657 when 733,
			1893043 when 734,
			1894425 when 735,
			1895803 when 736,
			1897176 when 737,
			1898545 when 738,
			1899909 when 739,
			1901269 when 740,
			1902624 when 741,
			1903975 when 742,
			1905322 when 743,
			1906663 when 744,
			1908001 when 745,
			1909334 when 746,
			1910662 when 747,
			1911986 when 748,
			1913306 when 749,
			1914620 when 750,
			1915931 when 751,
			1917237 when 752,
			1918538 when 753,
			1919835 when 754,
			1921127 when 755,
			1922415 when 756,
			1923699 when 757,
			1924977 when 758,
			1926252 when 759,
			1927521 when 760,
			1928787 when 761,
			1930047 when 762,
			1931303 when 763,
			1932555 when 764,
			1933802 when 765,
			1935045 when 766,
			1936282 when 767,
			1937516 when 768,
			1938745 when 769,
			1939969 when 770,
			1941189 when 771,
			1942404 when 772,
			1943614 when 773,
			1944820 when 774,
			1946022 when 775,
			1947218 when 776,
			1948411 when 777,
			1949598 when 778,
			1950781 when 779,
			1951960 when 780,
			1953134 when 781,
			1954303 when 782,
			1955468 when 783,
			1956628 when 784,
			1957783 when 785,
			1958934 when 786,
			1960080 when 787,
			1961222 when 788,
			1962359 when 789,
			1963491 when 790,
			1964619 when 791,
			1965742 when 792,
			1966861 when 793,
			1967975 when 794,
			1969084 when 795,
			1970189 when 796,
			1971289 when 797,
			1972384 when 798,
			1973475 when 799,
			1974561 when 800,
			1975642 when 801,
			1976719 when 802,
			1977791 when 803,
			1978859 when 804,
			1979922 when 805,
			1980980 when 806,
			1982033 when 807,
			1983082 when 808,
			1984126 when 809,
			1985166 when 810,
			1986201 when 811,
			1987231 when 812,
			1988257 when 813,
			1989277 when 814,
			1990293 when 815,
			1991305 when 816,
			1992312 when 817,
			1993314 when 818,
			1994311 when 819,
			1995304 when 820,
			1996292 when 821,
			1997275 when 822,
			1998254 when 823,
			1999228 when 824,
			2000197 when 825,
			2001161 when 826,
			2002121 when 827,
			2003076 when 828,
			2004027 when 829,
			2004972 when 830,
			2005913 when 831,
			2006849 when 832,
			2007781 when 833,
			2008708 when 834,
			2009630 when 835,
			2010547 when 836,
			2011459 when 837,
			2012367 when 838,
			2013270 when 839,
			2014169 when 840,
			2015062 when 841,
			2015951 when 842,
			2016835 when 843,
			2017715 when 844,
			2018589 when 845,
			2019459 when 846,
			2020325 when 847,
			2021185 when 848,
			2022041 when 849,
			2022891 when 850,
			2023738 when 851,
			2024579 when 852,
			2025415 when 853,
			2026247 when 854,
			2027074 when 855,
			2027897 when 856,
			2028714 when 857,
			2029527 when 858,
			2030335 when 859,
			2031138 when 860,
			2031936 when 861,
			2032730 when 862,
			2033519 when 863,
			2034303 when 864,
			2035082 when 865,
			2035857 when 866,
			2036626 when 867,
			2037391 when 868,
			2038151 when 869,
			2038907 when 870,
			2039657 when 871,
			2040403 when 872,
			2041144 when 873,
			2041880 when 874,
			2042611 when 875,
			2043338 when 876,
			2044059 when 877,
			2044776 when 878,
			2045488 when 879,
			2046196 when 880,
			2046898 when 881,
			2047596 when 882,
			2048289 when 883,
			2048977 when 884,
			2049660 when 885,
			2050338 when 886,
			2051012 when 887,
			2051680 when 888,
			2052344 when 889,
			2053003 when 890,
			2053657 when 891,
			2054307 when 892,
			2054951 when 893,
			2055591 when 894,
			2056226 when 895,
			2056856 when 896,
			2057481 when 897,
			2058101 when 898,
			2058717 when 899,
			2059327 when 900,
			2059933 when 901,
			2060534 when 902,
			2061130 when 903,
			2061722 when 904,
			2062308 when 905,
			2062890 when 906,
			2063466 when 907,
			2064038 when 908,
			2064605 when 909,
			2065167 when 910,
			2065725 when 911,
			2066277 when 912,
			2066825 when 913,
			2067367 when 914,
			2067905 when 915,
			2068438 when 916,
			2068966 when 917,
			2069489 when 918,
			2070008 when 919,
			2070521 when 920,
			2071030 when 921,
			2071533 when 922,
			2072032 when 923,
			2072526 when 924,
			2073015 when 925,
			2073500 when 926,
			2073979 when 927,
			2074453 when 928,
			2074923 when 929,
			2075388 when 930,
			2075848 when 931,
			2076303 when 932,
			2076753 when 933,
			2077198 when 934,
			2077638 when 935,
			2078073 when 936,
			2078504 when 937,
			2078930 when 938,
			2079350 when 939,
			2079766 when 940,
			2080177 when 941,
			2080583 when 942,
			2080984 when 943,
			2081380 when 944,
			2081772 when 945,
			2082158 when 946,
			2082540 when 947,
			2082916 when 948,
			2083288 when 949,
			2083655 when 950,
			2084017 when 951,
			2084374 when 952,
			2084726 when 953,
			2085073 when 954,
			2085416 when 955,
			2085753 when 956,
			2086086 when 957,
			2086413 when 958,
			2086736 when 959,
			2087054 when 960,
			2087367 when 961,
			2087674 when 962,
			2087977 when 963,
			2088276 when 964,
			2088569 when 965,
			2088857 when 966,
			2089141 when 967,
			2089419 when 968,
			2089693 when 969,
			2089961 when 970,
			2090225 when 971,
			2090484 when 972,
			2090738 when 973,
			2090987 when 974,
			2091231 when 975,
			2091470 when 976,
			2091704 when 977,
			2091933 when 978,
			2092157 when 979,
			2092377 when 980,
			2092591 when 981,
			2092801 when 982,
			2093006 when 983,
			2093205 when 984,
			2093400 when 985,
			2093590 when 986,
			2093775 when 987,
			2093955 when 988,
			2094130 when 989,
			2094300 when 990,
			2094466 when 991,
			2094626 when 992,
			2094781 when 993,
			2094932 when 994,
			2095077 when 995,
			2095218 when 996,
			2095354 when 997,
			2095484 when 998,
			2095610 when 999,
			2095731 when 1000,
			2095847 when 1001,
			2095958 when 1002,
			2096064 when 1003,
			2096165 when 1004,
			2096261 when 1005,
			2096353 when 1006,
			2096439 when 1007,
			2096520 when 1008,
			2096597 when 1009,
			2096668 when 1010,
			2096735 when 1011,
			2096797 when 1012,
			2096853 when 1013,
			2096905 when 1014,
			2096952 when 1015,
			2096994 when 1016,
			2097031 when 1017,
			2097063 when 1018,
			2097090 when 1019,
			2097113 when 1020,
			2097130 when 1021,
			2097142 when 1022,
			2097150 when 1023,
			2097152 when 1024,
			2097150 when 1025,
			2097142 when 1026,
			2097130 when 1027,
			2097113 when 1028,
			2097090 when 1029,
			2097063 when 1030,
			2097031 when 1031,
			2096994 when 1032,
			2096952 when 1033,
			2096905 when 1034,
			2096853 when 1035,
			2096797 when 1036,
			2096735 when 1037,
			2096668 when 1038,
			2096597 when 1039,
			2096520 when 1040,
			2096439 when 1041,
			2096353 when 1042,
			2096261 when 1043,
			2096165 when 1044,
			2096064 when 1045,
			2095958 when 1046,
			2095847 when 1047,
			2095731 when 1048,
			2095610 when 1049,
			2095484 when 1050,
			2095354 when 1051,
			2095218 when 1052,
			2095077 when 1053,
			2094932 when 1054,
			2094781 when 1055,
			2094626 when 1056,
			2094466 when 1057,
			2094300 when 1058,
			2094130 when 1059,
			2093955 when 1060,
			2093775 when 1061,
			2093590 when 1062,
			2093400 when 1063,
			2093205 when 1064,
			2093006 when 1065,
			2092801 when 1066,
			2092591 when 1067,
			2092377 when 1068,
			2092157 when 1069,
			2091933 when 1070,
			2091704 when 1071,
			2091470 when 1072,
			2091231 when 1073,
			2090987 when 1074,
			2090738 when 1075,
			2090484 when 1076,
			2090225 when 1077,
			2089961 when 1078,
			2089693 when 1079,
			2089419 when 1080,
			2089141 when 1081,
			2088857 when 1082,
			2088569 when 1083,
			2088276 when 1084,
			2087977 when 1085,
			2087674 when 1086,
			2087367 when 1087,
			2087054 when 1088,
			2086736 when 1089,
			2086413 when 1090,
			2086086 when 1091,
			2085753 when 1092,
			2085416 when 1093,
			2085073 when 1094,
			2084726 when 1095,
			2084374 when 1096,
			2084017 when 1097,
			2083655 when 1098,
			2083288 when 1099,
			2082916 when 1100,
			2082540 when 1101,
			2082158 when 1102,
			2081772 when 1103,
			2081380 when 1104,
			2080984 when 1105,
			2080583 when 1106,
			2080177 when 1107,
			2079766 when 1108,
			2079350 when 1109,
			2078930 when 1110,
			2078504 when 1111,
			2078073 when 1112,
			2077638 when 1113,
			2077198 when 1114,
			2076753 when 1115,
			2076303 when 1116,
			2075848 when 1117,
			2075388 when 1118,
			2074923 when 1119,
			2074453 when 1120,
			2073979 when 1121,
			2073500 when 1122,
			2073015 when 1123,
			2072526 when 1124,
			2072032 when 1125,
			2071533 when 1126,
			2071030 when 1127,
			2070521 when 1128,
			2070008 when 1129,
			2069489 when 1130,
			2068966 when 1131,
			2068438 when 1132,
			2067905 when 1133,
			2067367 when 1134,
			2066825 when 1135,
			2066277 when 1136,
			2065725 when 1137,
			2065167 when 1138,
			2064605 when 1139,
			2064038 when 1140,
			2063466 when 1141,
			2062890 when 1142,
			2062308 when 1143,
			2061722 when 1144,
			2061130 when 1145,
			2060534 when 1146,
			2059933 when 1147,
			2059327 when 1148,
			2058717 when 1149,
			2058101 when 1150,
			2057481 when 1151,
			2056856 when 1152,
			2056226 when 1153,
			2055591 when 1154,
			2054951 when 1155,
			2054307 when 1156,
			2053657 when 1157,
			2053003 when 1158,
			2052344 when 1159,
			2051680 when 1160,
			2051012 when 1161,
			2050338 when 1162,
			2049660 when 1163,
			2048977 when 1164,
			2048289 when 1165,
			2047596 when 1166,
			2046898 when 1167,
			2046196 when 1168,
			2045488 when 1169,
			2044776 when 1170,
			2044059 when 1171,
			2043338 when 1172,
			2042611 when 1173,
			2041880 when 1174,
			2041144 when 1175,
			2040403 when 1176,
			2039657 when 1177,
			2038907 when 1178,
			2038151 when 1179,
			2037391 when 1180,
			2036626 when 1181,
			2035857 when 1182,
			2035082 when 1183,
			2034303 when 1184,
			2033519 when 1185,
			2032730 when 1186,
			2031936 when 1187,
			2031138 when 1188,
			2030335 when 1189,
			2029527 when 1190,
			2028714 when 1191,
			2027897 when 1192,
			2027074 when 1193,
			2026247 when 1194,
			2025415 when 1195,
			2024579 when 1196,
			2023738 when 1197,
			2022891 when 1198,
			2022041 when 1199,
			2021185 when 1200,
			2020325 when 1201,
			2019459 when 1202,
			2018589 when 1203,
			2017715 when 1204,
			2016835 when 1205,
			2015951 when 1206,
			2015062 when 1207,
			2014169 when 1208,
			2013270 when 1209,
			2012367 when 1210,
			2011459 when 1211,
			2010547 when 1212,
			2009630 when 1213,
			2008708 when 1214,
			2007781 when 1215,
			2006849 when 1216,
			2005913 when 1217,
			2004972 when 1218,
			2004027 when 1219,
			2003076 when 1220,
			2002121 when 1221,
			2001161 when 1222,
			2000197 when 1223,
			1999228 when 1224,
			1998254 when 1225,
			1997275 when 1226,
			1996292 when 1227,
			1995304 when 1228,
			1994311 when 1229,
			1993314 when 1230,
			1992312 when 1231,
			1991305 when 1232,
			1990293 when 1233,
			1989277 when 1234,
			1988257 when 1235,
			1987231 when 1236,
			1986201 when 1237,
			1985166 when 1238,
			1984126 when 1239,
			1983082 when 1240,
			1982033 when 1241,
			1980980 when 1242,
			1979922 when 1243,
			1978859 when 1244,
			1977791 when 1245,
			1976719 when 1246,
			1975642 when 1247,
			1974561 when 1248,
			1973475 when 1249,
			1972384 when 1250,
			1971289 when 1251,
			1970189 when 1252,
			1969084 when 1253,
			1967975 when 1254,
			1966861 when 1255,
			1965742 when 1256,
			1964619 when 1257,
			1963491 when 1258,
			1962359 when 1259,
			1961222 when 1260,
			1960080 when 1261,
			1958934 when 1262,
			1957783 when 1263,
			1956628 when 1264,
			1955468 when 1265,
			1954303 when 1266,
			1953134 when 1267,
			1951960 when 1268,
			1950781 when 1269,
			1949598 when 1270,
			1948411 when 1271,
			1947218 when 1272,
			1946022 when 1273,
			1944820 when 1274,
			1943614 when 1275,
			1942404 when 1276,
			1941189 when 1277,
			1939969 when 1278,
			1938745 when 1279,
			1937516 when 1280,
			1936282 when 1281,
			1935045 when 1282,
			1933802 when 1283,
			1932555 when 1284,
			1931303 when 1285,
			1930047 when 1286,
			1928787 when 1287,
			1927521 when 1288,
			1926252 when 1289,
			1924977 when 1290,
			1923699 when 1291,
			1922415 when 1292,
			1921127 when 1293,
			1919835 when 1294,
			1918538 when 1295,
			1917237 when 1296,
			1915931 when 1297,
			1914620 when 1298,
			1913306 when 1299,
			1911986 when 1300,
			1910662 when 1301,
			1909334 when 1302,
			1908001 when 1303,
			1906663 when 1304,
			1905322 when 1305,
			1903975 when 1306,
			1902624 when 1307,
			1901269 when 1308,
			1899909 when 1309,
			1898545 when 1310,
			1897176 when 1311,
			1895803 when 1312,
			1894425 when 1313,
			1893043 when 1314,
			1891657 when 1315,
			1890266 when 1316,
			1888870 when 1317,
			1887470 when 1318,
			1886066 when 1319,
			1884657 when 1320,
			1883244 when 1321,
			1881826 when 1322,
			1880404 when 1323,
			1878977 when 1324,
			1877546 when 1325,
			1876111 when 1326,
			1874671 when 1327,
			1873227 when 1328,
			1871779 when 1329,
			1870326 when 1330,
			1868868 when 1331,
			1867406 when 1332,
			1865940 when 1333,
			1864470 when 1334,
			1862995 when 1335,
			1861515 when 1336,
			1860031 when 1337,
			1858543 when 1338,
			1857051 when 1339,
			1855554 when 1340,
			1854053 when 1341,
			1852547 when 1342,
			1851037 when 1343,
			1849523 when 1344,
			1848004 when 1345,
			1846481 when 1346,
			1844954 when 1347,
			1843422 when 1348,
			1841886 when 1349,
			1840346 when 1350,
			1838801 when 1351,
			1837252 when 1352,
			1835699 when 1353,
			1834141 when 1354,
			1832579 when 1355,
			1831013 when 1356,
			1829442 when 1357,
			1827867 when 1358,
			1826288 when 1359,
			1824705 when 1360,
			1823117 when 1361,
			1821525 when 1362,
			1819928 when 1363,
			1818328 when 1364,
			1816723 when 1365,
			1815114 when 1366,
			1813500 when 1367,
			1811882 when 1368,
			1810260 when 1369,
			1808634 when 1370,
			1807004 when 1371,
			1805369 when 1372,
			1803730 when 1373,
			1802087 when 1374,
			1800439 when 1375,
			1798787 when 1376,
			1797131 when 1377,
			1795471 when 1378,
			1793807 when 1379,
			1792138 when 1380,
			1790465 when 1381,
			1788788 when 1382,
			1787107 when 1383,
			1785421 when 1384,
			1783732 when 1385,
			1782038 when 1386,
			1780340 when 1387,
			1778637 when 1388,
			1776931 when 1389,
			1775220 when 1390,
			1773505 when 1391,
			1771786 when 1392,
			1770063 when 1393,
			1768336 when 1394,
			1766604 when 1395,
			1764869 when 1396,
			1763129 when 1397,
			1761385 when 1398,
			1759637 when 1399,
			1757885 when 1400,
			1756128 when 1401,
			1754368 when 1402,
			1752603 when 1403,
			1750834 when 1404,
			1749061 when 1405,
			1747284 when 1406,
			1745503 when 1407,
			1743718 when 1408,
			1741929 when 1409,
			1740135 when 1410,
			1738338 when 1411,
			1736536 when 1412,
			1734731 when 1413,
			1732921 when 1414,
			1731107 when 1415,
			1729289 when 1416,
			1727467 when 1417,
			1725641 when 1418,
			1723811 when 1419,
			1721977 when 1420,
			1720139 when 1421,
			1718296 when 1422,
			1716450 when 1423,
			1714600 when 1424,
			1712745 when 1425,
			1710887 when 1426,
			1709024 when 1427,
			1707158 when 1428,
			1705287 when 1429,
			1703413 when 1430,
			1701534 when 1431,
			1699652 when 1432,
			1697765 when 1433,
			1695875 when 1434,
			1693980 when 1435,
			1692082 when 1436,
			1690180 when 1437,
			1688273 when 1438,
			1686363 when 1439,
			1684448 when 1440,
			1682530 when 1441,
			1680608 when 1442,
			1678681 when 1443,
			1676751 when 1444,
			1674817 when 1445,
			1672879 when 1446,
			1670937 when 1447,
			1668991 when 1448,
			1667041 when 1449,
			1665087 when 1450,
			1663130 when 1451,
			1661168 when 1452,
			1659202 when 1453,
			1657233 when 1454,
			1655260 when 1455,
			1653282 when 1456,
			1651301 when 1457,
			1649316 when 1458,
			1647327 when 1459,
			1645334 when 1460,
			1643338 when 1461,
			1641337 when 1462,
			1639333 when 1463,
			1637325 when 1464,
			1635313 when 1465,
			1633297 when 1466,
			1631277 when 1467,
			1629253 when 1468,
			1627226 when 1469,
			1625194 when 1470,
			1623159 when 1471,
			1621120 when 1472,
			1619078 when 1473,
			1617031 when 1474,
			1614981 when 1475,
			1612927 when 1476,
			1610869 when 1477,
			1608807 when 1478,
			1606741 when 1479,
			1604672 when 1480,
			1602599 when 1481,
			1600522 when 1482,
			1598441 when 1483,
			1596357 when 1484,
			1594269 when 1485,
			1592177 when 1486,
			1590081 when 1487,
			1587982 when 1488,
			1585879 when 1489,
			1583772 when 1490,
			1581662 when 1491,
			1579547 when 1492,
			1577429 when 1493,
			1575307 when 1494,
			1573182 when 1495,
			1571053 when 1496,
			1568920 when 1497,
			1566784 when 1498,
			1564643 when 1499,
			1562499 when 1500,
			1560352 when 1501,
			1558201 when 1502,
			1556046 when 1503,
			1553887 when 1504,
			1551725 when 1505,
			1549559 when 1506,
			1547390 when 1507,
			1545216 when 1508,
			1543040 when 1509,
			1540859 when 1510,
			1538675 when 1511,
			1536487 when 1512,
			1534296 when 1513,
			1532101 when 1514,
			1529903 when 1515,
			1527701 when 1516,
			1525495 when 1517,
			1523286 when 1518,
			1521073 when 1519,
			1518856 when 1520,
			1516636 when 1521,
			1514413 when 1522,
			1512185 when 1523,
			1509955 when 1524,
			1507720 when 1525,
			1505483 when 1526,
			1503241 when 1527,
			1500996 when 1528,
			1498748 when 1529,
			1496496 when 1530,
			1494240 when 1531,
			1491981 when 1532,
			1489719 when 1533,
			1487453 when 1534,
			1485183 when 1535,
			1482910 when 1536,
			1480634 when 1537,
			1478354 when 1538,
			1476070 when 1539,
			1473784 when 1540,
			1471493 when 1541,
			1469199 when 1542,
			1466902 when 1543,
			1464601 when 1544,
			1462297 when 1545,
			1459989 when 1546,
			1457678 when 1547,
			1455364 when 1548,
			1453046 when 1549,
			1450724 when 1550,
			1448400 when 1551,
			1446071 when 1552,
			1443740 when 1553,
			1441405 when 1554,
			1439066 when 1555,
			1436725 when 1556,
			1434379 when 1557,
			1432031 when 1558,
			1429679 when 1559,
			1427324 when 1560,
			1424965 when 1561,
			1422603 when 1562,
			1420238 when 1563,
			1417869 when 1564,
			1415497 when 1565,
			1413122 when 1566,
			1410743 when 1567,
			1408361 when 1568,
			1405976 when 1569,
			1403587 when 1570,
			1401195 when 1571,
			1398800 when 1572,
			1396402 when 1573,
			1394000 when 1574,
			1391595 when 1575,
			1389187 when 1576,
			1386775 when 1577,
			1384360 when 1578,
			1381942 when 1579,
			1379521 when 1580,
			1377096 when 1581,
			1374668 when 1582,
			1372237 when 1583,
			1369803 when 1584,
			1367365 when 1585,
			1364924 when 1586,
			1362480 when 1587,
			1360033 when 1588,
			1357583 when 1589,
			1355129 when 1590,
			1352673 when 1591,
			1350213 when 1592,
			1347749 when 1593,
			1345283 when 1594,
			1342814 when 1595,
			1340341 when 1596,
			1337865 when 1597,
			1335386 when 1598,
			1332904 when 1599,
			1330419 when 1600,
			1327931 when 1601,
			1325439 when 1602,
			1322945 when 1603,
			1320447 when 1604,
			1317946 when 1605,
			1315442 when 1606,
			1312935 when 1607,
			1310425 when 1608,
			1307912 when 1609,
			1305396 when 1610,
			1302877 when 1611,
			1300354 when 1612,
			1297829 when 1613,
			1295300 when 1614,
			1292769 when 1615,
			1290234 when 1616,
			1287697 when 1617,
			1285156 when 1618,
			1282612 when 1619,
			1280066 when 1620,
			1277516 when 1621,
			1274963 when 1622,
			1272407 when 1623,
			1269849 when 1624,
			1267287 when 1625,
			1264722 when 1626,
			1262155 when 1627,
			1259584 when 1628,
			1257010 when 1629,
			1254434 when 1630,
			1251854 when 1631,
			1249272 when 1632,
			1246687 when 1633,
			1244098 when 1634,
			1241507 when 1635,
			1238913 when 1636,
			1236316 when 1637,
			1233716 when 1638,
			1231113 when 1639,
			1228507 when 1640,
			1225898 when 1641,
			1223287 when 1642,
			1220672 when 1643,
			1218055 when 1644,
			1215435 when 1645,
			1212812 when 1646,
			1210186 when 1647,
			1207557 when 1648,
			1204926 when 1649,
			1202291 when 1650,
			1199654 when 1651,
			1197014 when 1652,
			1194371 when 1653,
			1191725 when 1654,
			1189077 when 1655,
			1186426 when 1656,
			1183772 when 1657,
			1181115 when 1658,
			1178455 when 1659,
			1175793 when 1660,
			1173127 when 1661,
			1170459 when 1662,
			1167789 when 1663,
			1165115 when 1664,
			1162439 when 1665,
			1159760 when 1666,
			1157078 when 1667,
			1154394 when 1668,
			1151707 when 1669,
			1149017 when 1670,
			1146325 when 1671,
			1143629 when 1672,
			1140931 when 1673,
			1138231 when 1674,
			1135528 when 1675,
			1132822 when 1676,
			1130113 when 1677,
			1127402 when 1678,
			1124688 when 1679,
			1121971 when 1680,
			1119252 when 1681,
			1116530 when 1682,
			1113806 when 1683,
			1111079 when 1684,
			1108349 when 1685,
			1105617 when 1686,
			1102882 when 1687,
			1100144 when 1688,
			1097404 when 1689,
			1094662 when 1690,
			1091916 when 1691,
			1089168 when 1692,
			1086418 when 1693,
			1083665 when 1694,
			1080910 when 1695,
			1078152 when 1696,
			1075391 when 1697,
			1072628 when 1698,
			1069862 when 1699,
			1067094 when 1700,
			1064323 when 1701,
			1061550 when 1702,
			1058775 when 1703,
			1055997 when 1704,
			1053216 when 1705,
			1050433 when 1706,
			1047647 when 1707,
			1044859 when 1708,
			1042069 when 1709,
			1039276 when 1710,
			1036480 when 1711,
			1033682 when 1712,
			1030882 when 1713,
			1028079 when 1714,
			1025274 when 1715,
			1022467 when 1716,
			1019657 when 1717,
			1016845 when 1718,
			1014030 when 1719,
			1011213 when 1720,
			1008393 when 1721,
			1005571 when 1722,
			1002747 when 1723,
			999920 when 1724,
			997092 when 1725,
			994260 when 1726,
			991427 when 1727,
			988591 when 1728,
			985752 when 1729,
			982912 when 1730,
			980069 when 1731,
			977224 when 1732,
			974376 when 1733,
			971526 when 1734,
			968674 when 1735,
			965820 when 1736,
			962963 when 1737,
			960104 when 1738,
			957243 when 1739,
			954379 when 1740,
			951514 when 1741,
			948646 when 1742,
			945776 when 1743,
			942903 when 1744,
			940029 when 1745,
			937152 when 1746,
			934273 when 1747,
			931392 when 1748,
			928508 when 1749,
			925623 when 1750,
			922735 when 1751,
			919845 when 1752,
			916953 when 1753,
			914059 when 1754,
			911162 when 1755,
			908264 when 1756,
			905363 when 1757,
			902460 when 1758,
			899555 when 1759,
			896648 when 1760,
			893739 when 1761,
			890828 when 1762,
			887914 when 1763,
			884999 when 1764,
			882081 when 1765,
			879162 when 1766,
			876240 when 1767,
			873316 when 1768,
			870390 when 1769,
			867462 when 1770,
			864533 when 1771,
			861601 when 1772,
			858667 when 1773,
			855731 when 1774,
			852793 when 1775,
			849853 when 1776,
			846911 when 1777,
			843967 when 1778,
			841021 when 1779,
			838073 when 1780,
			835123 when 1781,
			832171 when 1782,
			829217 when 1783,
			826261 when 1784,
			823303 when 1785,
			820344 when 1786,
			817382 when 1787,
			814419 when 1788,
			811453 when 1789,
			808486 when 1790,
			805516 when 1791,
			802545 when 1792,
			799572 when 1793,
			796597 when 1794,
			793621 when 1795,
			790642 when 1796,
			787661 when 1797,
			784679 when 1798,
			781695 when 1799,
			778709 when 1800,
			775721 when 1801,
			772731 when 1802,
			769739 when 1803,
			766746 when 1804,
			763751 when 1805,
			760754 when 1806,
			757755 when 1807,
			754755 when 1808,
			751752 when 1809,
			748748 when 1810,
			745742 when 1811,
			742735 when 1812,
			739725 when 1813,
			736714 when 1814,
			733701 when 1815,
			730687 when 1816,
			727671 when 1817,
			724653 when 1818,
			721633 when 1819,
			718612 when 1820,
			715589 when 1821,
			712564 when 1822,
			709537 when 1823,
			706509 when 1824,
			703479 when 1825,
			700448 when 1826,
			697415 when 1827,
			694380 when 1828,
			691344 when 1829,
			688306 when 1830,
			685266 when 1831,
			682225 when 1832,
			679182 when 1833,
			676138 when 1834,
			673092 when 1835,
			670044 when 1836,
			666995 when 1837,
			663944 when 1838,
			660892 when 1839,
			657838 when 1840,
			654783 when 1841,
			651726 when 1842,
			648667 when 1843,
			645607 when 1844,
			642546 when 1845,
			639483 when 1846,
			636418 when 1847,
			633352 when 1848,
			630285 when 1849,
			627216 when 1850,
			624145 when 1851,
			621073 when 1852,
			618000 when 1853,
			614925 when 1854,
			611849 when 1855,
			608771 when 1856,
			605692 when 1857,
			602611 when 1858,
			599529 when 1859,
			596446 when 1860,
			593361 when 1861,
			590275 when 1862,
			587187 when 1863,
			584098 when 1864,
			581008 when 1865,
			577916 when 1866,
			574823 when 1867,
			571728 when 1868,
			568633 when 1869,
			565535 when 1870,
			562437 when 1871,
			559337 when 1872,
			556236 when 1873,
			553134 when 1874,
			550030 when 1875,
			546925 when 1876,
			543819 when 1877,
			540711 when 1878,
			537602 when 1879,
			534492 when 1880,
			531381 when 1881,
			528268 when 1882,
			525154 when 1883,
			522039 when 1884,
			518923 when 1885,
			515805 when 1886,
			512686 when 1887,
			509566 when 1888,
			506445 when 1889,
			503323 when 1890,
			500199 when 1891,
			497075 when 1892,
			493949 when 1893,
			490822 when 1894,
			487693 when 1895,
			484564 when 1896,
			481433 when 1897,
			478302 when 1898,
			475169 when 1899,
			472035 when 1900,
			468900 when 1901,
			465764 when 1902,
			462627 when 1903,
			459489 when 1904,
			456349 when 1905,
			453209 when 1906,
			450067 when 1907,
			446925 when 1908,
			443781 when 1909,
			440636 when 1910,
			437491 when 1911,
			434344 when 1912,
			431196 when 1913,
			428048 when 1914,
			424898 when 1915,
			421747 when 1916,
			418595 when 1917,
			415442 when 1918,
			412289 when 1919,
			409134 when 1920,
			405978 when 1921,
			402822 when 1922,
			399664 when 1923,
			396506 when 1924,
			393346 when 1925,
			390186 when 1926,
			387025 when 1927,
			383862 when 1928,
			380699 when 1929,
			377535 when 1930,
			374371 when 1931,
			371205 when 1932,
			368038 when 1933,
			364871 when 1934,
			361702 when 1935,
			358533 when 1936,
			355363 when 1937,
			352192 when 1938,
			349020 when 1939,
			345848 when 1940,
			342675 when 1941,
			339500 when 1942,
			336325 when 1943,
			333150 when 1944,
			329973 when 1945,
			326796 when 1946,
			323618 when 1947,
			320439 when 1948,
			317259 when 1949,
			314079 when 1950,
			310898 when 1951,
			307716 when 1952,
			304534 when 1953,
			301350 when 1954,
			298166 when 1955,
			294982 when 1956,
			291796 when 1957,
			288610 when 1958,
			285424 when 1959,
			282236 when 1960,
			279048 when 1961,
			275859 when 1962,
			272670 when 1963,
			269480 when 1964,
			266289 when 1965,
			263098 when 1966,
			259906 when 1967,
			256714 when 1968,
			253521 when 1969,
			250327 when 1970,
			247133 when 1971,
			243938 when 1972,
			240742 when 1973,
			237546 when 1974,
			234350 when 1975,
			231153 when 1976,
			227955 when 1977,
			224757 when 1978,
			221558 when 1979,
			218359 when 1980,
			215159 when 1981,
			211959 when 1982,
			208758 when 1983,
			205557 when 1984,
			202355 when 1985,
			199153 when 1986,
			195950 when 1987,
			192747 when 1988,
			189543 when 1989,
			186339 when 1990,
			183135 when 1991,
			179930 when 1992,
			176725 when 1993,
			173519 when 1994,
			170313 when 1995,
			167106 when 1996,
			163899 when 1997,
			160692 when 1998,
			157484 when 1999,
			154276 when 2000,
			151068 when 2001,
			147859 when 2002,
			144650 when 2003,
			141440 when 2004,
			138230 when 2005,
			135020 when 2006,
			131810 when 2007,
			128599 when 2008,
			125388 when 2009,
			122176 when 2010,
			118965 when 2011,
			115753 when 2012,
			112541 when 2013,
			109328 when 2014,
			106115 when 2015,
			102902 when 2016,
			99689 when 2017,
			96476 when 2018,
			93262 when 2019,
			90048 when 2020,
			86834 when 2021,
			83620 when 2022,
			80405 when 2023,
			77190 when 2024,
			73975 when 2025,
			70760 when 2026,
			67545 when 2027,
			64330 when 2028,
			61114 when 2029,
			57898 when 2030,
			54683 when 2031,
			51467 when 2032,
			48251 when 2033,
			45034 when 2034,
			41818 when 2035,
			38602 when 2036,
			35385 when 2037,
			32169 when 2038,
			28952 when 2039,
			25735 when 2040,
			22519 when 2041,
			19302 when 2042,
			16085 when 2043,
			12868 when 2044,
			9651 when 2045,
			6434 when 2046,
			3217 when 2047,
			0 when 2048,
			-3217 when 2049,
			-6434 when 2050,
			-9651 when 2051,
			-12868 when 2052,
			-16085 when 2053,
			-19302 when 2054,
			-22519 when 2055,
			-25735 when 2056,
			-28952 when 2057,
			-32169 when 2058,
			-35385 when 2059,
			-38602 when 2060,
			-41818 when 2061,
			-45034 when 2062,
			-48251 when 2063,
			-51467 when 2064,
			-54683 when 2065,
			-57898 when 2066,
			-61114 when 2067,
			-64330 when 2068,
			-67545 when 2069,
			-70760 when 2070,
			-73975 when 2071,
			-77190 when 2072,
			-80405 when 2073,
			-83620 when 2074,
			-86834 when 2075,
			-90048 when 2076,
			-93262 when 2077,
			-96476 when 2078,
			-99689 when 2079,
			-102902 when 2080,
			-106115 when 2081,
			-109328 when 2082,
			-112541 when 2083,
			-115753 when 2084,
			-118965 when 2085,
			-122176 when 2086,
			-125388 when 2087,
			-128599 when 2088,
			-131810 when 2089,
			-135020 when 2090,
			-138230 when 2091,
			-141440 when 2092,
			-144650 when 2093,
			-147859 when 2094,
			-151068 when 2095,
			-154276 when 2096,
			-157484 when 2097,
			-160692 when 2098,
			-163899 when 2099,
			-167106 when 2100,
			-170313 when 2101,
			-173519 when 2102,
			-176725 when 2103,
			-179930 when 2104,
			-183135 when 2105,
			-186339 when 2106,
			-189543 when 2107,
			-192747 when 2108,
			-195950 when 2109,
			-199153 when 2110,
			-202355 when 2111,
			-205557 when 2112,
			-208758 when 2113,
			-211959 when 2114,
			-215159 when 2115,
			-218359 when 2116,
			-221558 when 2117,
			-224757 when 2118,
			-227955 when 2119,
			-231153 when 2120,
			-234350 when 2121,
			-237546 when 2122,
			-240742 when 2123,
			-243938 when 2124,
			-247133 when 2125,
			-250327 when 2126,
			-253521 when 2127,
			-256714 when 2128,
			-259906 when 2129,
			-263098 when 2130,
			-266289 when 2131,
			-269480 when 2132,
			-272670 when 2133,
			-275859 when 2134,
			-279048 when 2135,
			-282236 when 2136,
			-285424 when 2137,
			-288610 when 2138,
			-291796 when 2139,
			-294982 when 2140,
			-298166 when 2141,
			-301350 when 2142,
			-304534 when 2143,
			-307716 when 2144,
			-310898 when 2145,
			-314079 when 2146,
			-317259 when 2147,
			-320439 when 2148,
			-323618 when 2149,
			-326796 when 2150,
			-329973 when 2151,
			-333150 when 2152,
			-336325 when 2153,
			-339500 when 2154,
			-342675 when 2155,
			-345848 when 2156,
			-349020 when 2157,
			-352192 when 2158,
			-355363 when 2159,
			-358533 when 2160,
			-361702 when 2161,
			-364871 when 2162,
			-368038 when 2163,
			-371205 when 2164,
			-374371 when 2165,
			-377535 when 2166,
			-380699 when 2167,
			-383862 when 2168,
			-387025 when 2169,
			-390186 when 2170,
			-393346 when 2171,
			-396506 when 2172,
			-399664 when 2173,
			-402822 when 2174,
			-405978 when 2175,
			-409134 when 2176,
			-412289 when 2177,
			-415442 when 2178,
			-418595 when 2179,
			-421747 when 2180,
			-424898 when 2181,
			-428048 when 2182,
			-431196 when 2183,
			-434344 when 2184,
			-437491 when 2185,
			-440636 when 2186,
			-443781 when 2187,
			-446925 when 2188,
			-450067 when 2189,
			-453209 when 2190,
			-456349 when 2191,
			-459489 when 2192,
			-462627 when 2193,
			-465764 when 2194,
			-468900 when 2195,
			-472035 when 2196,
			-475169 when 2197,
			-478302 when 2198,
			-481433 when 2199,
			-484564 when 2200,
			-487693 when 2201,
			-490822 when 2202,
			-493949 when 2203,
			-497075 when 2204,
			-500199 when 2205,
			-503323 when 2206,
			-506445 when 2207,
			-509566 when 2208,
			-512686 when 2209,
			-515805 when 2210,
			-518923 when 2211,
			-522039 when 2212,
			-525154 when 2213,
			-528268 when 2214,
			-531381 when 2215,
			-534492 when 2216,
			-537602 when 2217,
			-540711 when 2218,
			-543819 when 2219,
			-546925 when 2220,
			-550030 when 2221,
			-553134 when 2222,
			-556236 when 2223,
			-559337 when 2224,
			-562437 when 2225,
			-565535 when 2226,
			-568633 when 2227,
			-571728 when 2228,
			-574823 when 2229,
			-577916 when 2230,
			-581008 when 2231,
			-584098 when 2232,
			-587187 when 2233,
			-590275 when 2234,
			-593361 when 2235,
			-596446 when 2236,
			-599529 when 2237,
			-602611 when 2238,
			-605692 when 2239,
			-608771 when 2240,
			-611849 when 2241,
			-614925 when 2242,
			-618000 when 2243,
			-621073 when 2244,
			-624145 when 2245,
			-627216 when 2246,
			-630285 when 2247,
			-633352 when 2248,
			-636418 when 2249,
			-639483 when 2250,
			-642546 when 2251,
			-645607 when 2252,
			-648667 when 2253,
			-651726 when 2254,
			-654783 when 2255,
			-657838 when 2256,
			-660892 when 2257,
			-663944 when 2258,
			-666995 when 2259,
			-670044 when 2260,
			-673092 when 2261,
			-676138 when 2262,
			-679182 when 2263,
			-682225 when 2264,
			-685266 when 2265,
			-688306 when 2266,
			-691344 when 2267,
			-694380 when 2268,
			-697415 when 2269,
			-700448 when 2270,
			-703479 when 2271,
			-706509 when 2272,
			-709537 when 2273,
			-712564 when 2274,
			-715589 when 2275,
			-718612 when 2276,
			-721633 when 2277,
			-724653 when 2278,
			-727671 when 2279,
			-730687 when 2280,
			-733701 when 2281,
			-736714 when 2282,
			-739725 when 2283,
			-742735 when 2284,
			-745742 when 2285,
			-748748 when 2286,
			-751752 when 2287,
			-754755 when 2288,
			-757755 when 2289,
			-760754 when 2290,
			-763751 when 2291,
			-766746 when 2292,
			-769739 when 2293,
			-772731 when 2294,
			-775721 when 2295,
			-778709 when 2296,
			-781695 when 2297,
			-784679 when 2298,
			-787661 when 2299,
			-790642 when 2300,
			-793621 when 2301,
			-796597 when 2302,
			-799572 when 2303,
			-802545 when 2304,
			-805516 when 2305,
			-808486 when 2306,
			-811453 when 2307,
			-814419 when 2308,
			-817382 when 2309,
			-820344 when 2310,
			-823303 when 2311,
			-826261 when 2312,
			-829217 when 2313,
			-832171 when 2314,
			-835123 when 2315,
			-838073 when 2316,
			-841021 when 2317,
			-843967 when 2318,
			-846911 when 2319,
			-849853 when 2320,
			-852793 when 2321,
			-855731 when 2322,
			-858667 when 2323,
			-861601 when 2324,
			-864533 when 2325,
			-867462 when 2326,
			-870390 when 2327,
			-873316 when 2328,
			-876240 when 2329,
			-879162 when 2330,
			-882081 when 2331,
			-884999 when 2332,
			-887914 when 2333,
			-890828 when 2334,
			-893739 when 2335,
			-896648 when 2336,
			-899555 when 2337,
			-902460 when 2338,
			-905363 when 2339,
			-908264 when 2340,
			-911162 when 2341,
			-914059 when 2342,
			-916953 when 2343,
			-919845 when 2344,
			-922735 when 2345,
			-925623 when 2346,
			-928508 when 2347,
			-931392 when 2348,
			-934273 when 2349,
			-937152 when 2350,
			-940029 when 2351,
			-942903 when 2352,
			-945776 when 2353,
			-948646 when 2354,
			-951514 when 2355,
			-954379 when 2356,
			-957243 when 2357,
			-960104 when 2358,
			-962963 when 2359,
			-965820 when 2360,
			-968674 when 2361,
			-971526 when 2362,
			-974376 when 2363,
			-977224 when 2364,
			-980069 when 2365,
			-982912 when 2366,
			-985752 when 2367,
			-988591 when 2368,
			-991427 when 2369,
			-994260 when 2370,
			-997092 when 2371,
			-999920 when 2372,
			-1002747 when 2373,
			-1005571 when 2374,
			-1008393 when 2375,
			-1011213 when 2376,
			-1014030 when 2377,
			-1016845 when 2378,
			-1019657 when 2379,
			-1022467 when 2380,
			-1025274 when 2381,
			-1028079 when 2382,
			-1030882 when 2383,
			-1033682 when 2384,
			-1036480 when 2385,
			-1039276 when 2386,
			-1042069 when 2387,
			-1044859 when 2388,
			-1047647 when 2389,
			-1050433 when 2390,
			-1053216 when 2391,
			-1055997 when 2392,
			-1058775 when 2393,
			-1061550 when 2394,
			-1064323 when 2395,
			-1067094 when 2396,
			-1069862 when 2397,
			-1072628 when 2398,
			-1075391 when 2399,
			-1078152 when 2400,
			-1080910 when 2401,
			-1083665 when 2402,
			-1086418 when 2403,
			-1089168 when 2404,
			-1091916 when 2405,
			-1094662 when 2406,
			-1097404 when 2407,
			-1100144 when 2408,
			-1102882 when 2409,
			-1105617 when 2410,
			-1108349 when 2411,
			-1111079 when 2412,
			-1113806 when 2413,
			-1116530 when 2414,
			-1119252 when 2415,
			-1121971 when 2416,
			-1124688 when 2417,
			-1127402 when 2418,
			-1130113 when 2419,
			-1132822 when 2420,
			-1135528 when 2421,
			-1138231 when 2422,
			-1140931 when 2423,
			-1143629 when 2424,
			-1146325 when 2425,
			-1149017 when 2426,
			-1151707 when 2427,
			-1154394 when 2428,
			-1157078 when 2429,
			-1159760 when 2430,
			-1162439 when 2431,
			-1165115 when 2432,
			-1167789 when 2433,
			-1170459 when 2434,
			-1173127 when 2435,
			-1175793 when 2436,
			-1178455 when 2437,
			-1181115 when 2438,
			-1183772 when 2439,
			-1186426 when 2440,
			-1189077 when 2441,
			-1191725 when 2442,
			-1194371 when 2443,
			-1197014 when 2444,
			-1199654 when 2445,
			-1202291 when 2446,
			-1204926 when 2447,
			-1207557 when 2448,
			-1210186 when 2449,
			-1212812 when 2450,
			-1215435 when 2451,
			-1218055 when 2452,
			-1220672 when 2453,
			-1223287 when 2454,
			-1225898 when 2455,
			-1228507 when 2456,
			-1231113 when 2457,
			-1233716 when 2458,
			-1236316 when 2459,
			-1238913 when 2460,
			-1241507 when 2461,
			-1244098 when 2462,
			-1246687 when 2463,
			-1249272 when 2464,
			-1251854 when 2465,
			-1254434 when 2466,
			-1257010 when 2467,
			-1259584 when 2468,
			-1262155 when 2469,
			-1264722 when 2470,
			-1267287 when 2471,
			-1269849 when 2472,
			-1272407 when 2473,
			-1274963 when 2474,
			-1277516 when 2475,
			-1280066 when 2476,
			-1282612 when 2477,
			-1285156 when 2478,
			-1287697 when 2479,
			-1290234 when 2480,
			-1292769 when 2481,
			-1295300 when 2482,
			-1297829 when 2483,
			-1300354 when 2484,
			-1302877 when 2485,
			-1305396 when 2486,
			-1307912 when 2487,
			-1310425 when 2488,
			-1312935 when 2489,
			-1315442 when 2490,
			-1317946 when 2491,
			-1320447 when 2492,
			-1322945 when 2493,
			-1325439 when 2494,
			-1327931 when 2495,
			-1330419 when 2496,
			-1332904 when 2497,
			-1335386 when 2498,
			-1337865 when 2499,
			-1340341 when 2500,
			-1342814 when 2501,
			-1345283 when 2502,
			-1347749 when 2503,
			-1350213 when 2504,
			-1352673 when 2505,
			-1355129 when 2506,
			-1357583 when 2507,
			-1360033 when 2508,
			-1362480 when 2509,
			-1364924 when 2510,
			-1367365 when 2511,
			-1369803 when 2512,
			-1372237 when 2513,
			-1374668 when 2514,
			-1377096 when 2515,
			-1379521 when 2516,
			-1381942 when 2517,
			-1384360 when 2518,
			-1386775 when 2519,
			-1389187 when 2520,
			-1391595 when 2521,
			-1394000 when 2522,
			-1396402 when 2523,
			-1398800 when 2524,
			-1401195 when 2525,
			-1403587 when 2526,
			-1405976 when 2527,
			-1408361 when 2528,
			-1410743 when 2529,
			-1413122 when 2530,
			-1415497 when 2531,
			-1417869 when 2532,
			-1420238 when 2533,
			-1422603 when 2534,
			-1424965 when 2535,
			-1427324 when 2536,
			-1429679 when 2537,
			-1432031 when 2538,
			-1434379 when 2539,
			-1436725 when 2540,
			-1439066 when 2541,
			-1441405 when 2542,
			-1443740 when 2543,
			-1446071 when 2544,
			-1448400 when 2545,
			-1450724 when 2546,
			-1453046 when 2547,
			-1455364 when 2548,
			-1457678 when 2549,
			-1459989 when 2550,
			-1462297 when 2551,
			-1464601 when 2552,
			-1466902 when 2553,
			-1469199 when 2554,
			-1471493 when 2555,
			-1473784 when 2556,
			-1476070 when 2557,
			-1478354 when 2558,
			-1480634 when 2559,
			-1482910 when 2560,
			-1485183 when 2561,
			-1487453 when 2562,
			-1489719 when 2563,
			-1491981 when 2564,
			-1494240 when 2565,
			-1496496 when 2566,
			-1498748 when 2567,
			-1500996 when 2568,
			-1503241 when 2569,
			-1505483 when 2570,
			-1507720 when 2571,
			-1509955 when 2572,
			-1512185 when 2573,
			-1514413 when 2574,
			-1516636 when 2575,
			-1518856 when 2576,
			-1521073 when 2577,
			-1523286 when 2578,
			-1525495 when 2579,
			-1527701 when 2580,
			-1529903 when 2581,
			-1532101 when 2582,
			-1534296 when 2583,
			-1536487 when 2584,
			-1538675 when 2585,
			-1540859 when 2586,
			-1543040 when 2587,
			-1545216 when 2588,
			-1547390 when 2589,
			-1549559 when 2590,
			-1551725 when 2591,
			-1553887 when 2592,
			-1556046 when 2593,
			-1558201 when 2594,
			-1560352 when 2595,
			-1562499 when 2596,
			-1564643 when 2597,
			-1566784 when 2598,
			-1568920 when 2599,
			-1571053 when 2600,
			-1573182 when 2601,
			-1575307 when 2602,
			-1577429 when 2603,
			-1579547 when 2604,
			-1581662 when 2605,
			-1583772 when 2606,
			-1585879 when 2607,
			-1587982 when 2608,
			-1590081 when 2609,
			-1592177 when 2610,
			-1594269 when 2611,
			-1596357 when 2612,
			-1598441 when 2613,
			-1600522 when 2614,
			-1602599 when 2615,
			-1604672 when 2616,
			-1606741 when 2617,
			-1608807 when 2618,
			-1610869 when 2619,
			-1612927 when 2620,
			-1614981 when 2621,
			-1617031 when 2622,
			-1619078 when 2623,
			-1621120 when 2624,
			-1623159 when 2625,
			-1625194 when 2626,
			-1627226 when 2627,
			-1629253 when 2628,
			-1631277 when 2629,
			-1633297 when 2630,
			-1635313 when 2631,
			-1637325 when 2632,
			-1639333 when 2633,
			-1641337 when 2634,
			-1643338 when 2635,
			-1645334 when 2636,
			-1647327 when 2637,
			-1649316 when 2638,
			-1651301 when 2639,
			-1653282 when 2640,
			-1655260 when 2641,
			-1657233 when 2642,
			-1659202 when 2643,
			-1661168 when 2644,
			-1663130 when 2645,
			-1665087 when 2646,
			-1667041 when 2647,
			-1668991 when 2648,
			-1670937 when 2649,
			-1672879 when 2650,
			-1674817 when 2651,
			-1676751 when 2652,
			-1678681 when 2653,
			-1680608 when 2654,
			-1682530 when 2655,
			-1684448 when 2656,
			-1686363 when 2657,
			-1688273 when 2658,
			-1690180 when 2659,
			-1692082 when 2660,
			-1693980 when 2661,
			-1695875 when 2662,
			-1697765 when 2663,
			-1699652 when 2664,
			-1701534 when 2665,
			-1703413 when 2666,
			-1705287 when 2667,
			-1707158 when 2668,
			-1709024 when 2669,
			-1710887 when 2670,
			-1712745 when 2671,
			-1714600 when 2672,
			-1716450 when 2673,
			-1718296 when 2674,
			-1720139 when 2675,
			-1721977 when 2676,
			-1723811 when 2677,
			-1725641 when 2678,
			-1727467 when 2679,
			-1729289 when 2680,
			-1731107 when 2681,
			-1732921 when 2682,
			-1734731 when 2683,
			-1736536 when 2684,
			-1738338 when 2685,
			-1740135 when 2686,
			-1741929 when 2687,
			-1743718 when 2688,
			-1745503 when 2689,
			-1747284 when 2690,
			-1749061 when 2691,
			-1750834 when 2692,
			-1752603 when 2693,
			-1754368 when 2694,
			-1756128 when 2695,
			-1757885 when 2696,
			-1759637 when 2697,
			-1761385 when 2698,
			-1763129 when 2699,
			-1764869 when 2700,
			-1766604 when 2701,
			-1768336 when 2702,
			-1770063 when 2703,
			-1771786 when 2704,
			-1773505 when 2705,
			-1775220 when 2706,
			-1776931 when 2707,
			-1778637 when 2708,
			-1780340 when 2709,
			-1782038 when 2710,
			-1783732 when 2711,
			-1785421 when 2712,
			-1787107 when 2713,
			-1788788 when 2714,
			-1790465 when 2715,
			-1792138 when 2716,
			-1793807 when 2717,
			-1795471 when 2718,
			-1797131 when 2719,
			-1798787 when 2720,
			-1800439 when 2721,
			-1802087 when 2722,
			-1803730 when 2723,
			-1805369 when 2724,
			-1807004 when 2725,
			-1808634 when 2726,
			-1810260 when 2727,
			-1811882 when 2728,
			-1813500 when 2729,
			-1815114 when 2730,
			-1816723 when 2731,
			-1818328 when 2732,
			-1819928 when 2733,
			-1821525 when 2734,
			-1823117 when 2735,
			-1824705 when 2736,
			-1826288 when 2737,
			-1827867 when 2738,
			-1829442 when 2739,
			-1831013 when 2740,
			-1832579 when 2741,
			-1834141 when 2742,
			-1835699 when 2743,
			-1837252 when 2744,
			-1838801 when 2745,
			-1840346 when 2746,
			-1841886 when 2747,
			-1843422 when 2748,
			-1844954 when 2749,
			-1846481 when 2750,
			-1848004 when 2751,
			-1849523 when 2752,
			-1851037 when 2753,
			-1852547 when 2754,
			-1854053 when 2755,
			-1855554 when 2756,
			-1857051 when 2757,
			-1858543 when 2758,
			-1860031 when 2759,
			-1861515 when 2760,
			-1862995 when 2761,
			-1864470 when 2762,
			-1865940 when 2763,
			-1867406 when 2764,
			-1868868 when 2765,
			-1870326 when 2766,
			-1871779 when 2767,
			-1873227 when 2768,
			-1874671 when 2769,
			-1876111 when 2770,
			-1877546 when 2771,
			-1878977 when 2772,
			-1880404 when 2773,
			-1881826 when 2774,
			-1883244 when 2775,
			-1884657 when 2776,
			-1886066 when 2777,
			-1887470 when 2778,
			-1888870 when 2779,
			-1890266 when 2780,
			-1891657 when 2781,
			-1893043 when 2782,
			-1894425 when 2783,
			-1895803 when 2784,
			-1897176 when 2785,
			-1898545 when 2786,
			-1899909 when 2787,
			-1901269 when 2788,
			-1902624 when 2789,
			-1903975 when 2790,
			-1905322 when 2791,
			-1906663 when 2792,
			-1908001 when 2793,
			-1909334 when 2794,
			-1910662 when 2795,
			-1911986 when 2796,
			-1913306 when 2797,
			-1914620 when 2798,
			-1915931 when 2799,
			-1917237 when 2800,
			-1918538 when 2801,
			-1919835 when 2802,
			-1921127 when 2803,
			-1922415 when 2804,
			-1923699 when 2805,
			-1924977 when 2806,
			-1926252 when 2807,
			-1927521 when 2808,
			-1928787 when 2809,
			-1930047 when 2810,
			-1931303 when 2811,
			-1932555 when 2812,
			-1933802 when 2813,
			-1935045 when 2814,
			-1936282 when 2815,
			-1937516 when 2816,
			-1938745 when 2817,
			-1939969 when 2818,
			-1941189 when 2819,
			-1942404 when 2820,
			-1943614 when 2821,
			-1944820 when 2822,
			-1946022 when 2823,
			-1947218 when 2824,
			-1948411 when 2825,
			-1949598 when 2826,
			-1950781 when 2827,
			-1951960 when 2828,
			-1953134 when 2829,
			-1954303 when 2830,
			-1955468 when 2831,
			-1956628 when 2832,
			-1957783 when 2833,
			-1958934 when 2834,
			-1960080 when 2835,
			-1961222 when 2836,
			-1962359 when 2837,
			-1963491 when 2838,
			-1964619 when 2839,
			-1965742 when 2840,
			-1966861 when 2841,
			-1967975 when 2842,
			-1969084 when 2843,
			-1970189 when 2844,
			-1971289 when 2845,
			-1972384 when 2846,
			-1973475 when 2847,
			-1974561 when 2848,
			-1975642 when 2849,
			-1976719 when 2850,
			-1977791 when 2851,
			-1978859 when 2852,
			-1979922 when 2853,
			-1980980 when 2854,
			-1982033 when 2855,
			-1983082 when 2856,
			-1984126 when 2857,
			-1985166 when 2858,
			-1986201 when 2859,
			-1987231 when 2860,
			-1988257 when 2861,
			-1989277 when 2862,
			-1990293 when 2863,
			-1991305 when 2864,
			-1992312 when 2865,
			-1993314 when 2866,
			-1994311 when 2867,
			-1995304 when 2868,
			-1996292 when 2869,
			-1997275 when 2870,
			-1998254 when 2871,
			-1999228 when 2872,
			-2000197 when 2873,
			-2001161 when 2874,
			-2002121 when 2875,
			-2003076 when 2876,
			-2004027 when 2877,
			-2004972 when 2878,
			-2005913 when 2879,
			-2006849 when 2880,
			-2007781 when 2881,
			-2008708 when 2882,
			-2009630 when 2883,
			-2010547 when 2884,
			-2011459 when 2885,
			-2012367 when 2886,
			-2013270 when 2887,
			-2014169 when 2888,
			-2015062 when 2889,
			-2015951 when 2890,
			-2016835 when 2891,
			-2017715 when 2892,
			-2018589 when 2893,
			-2019459 when 2894,
			-2020325 when 2895,
			-2021185 when 2896,
			-2022041 when 2897,
			-2022891 when 2898,
			-2023738 when 2899,
			-2024579 when 2900,
			-2025415 when 2901,
			-2026247 when 2902,
			-2027074 when 2903,
			-2027897 when 2904,
			-2028714 when 2905,
			-2029527 when 2906,
			-2030335 when 2907,
			-2031138 when 2908,
			-2031936 when 2909,
			-2032730 when 2910,
			-2033519 when 2911,
			-2034303 when 2912,
			-2035082 when 2913,
			-2035857 when 2914,
			-2036626 when 2915,
			-2037391 when 2916,
			-2038151 when 2917,
			-2038907 when 2918,
			-2039657 when 2919,
			-2040403 when 2920,
			-2041144 when 2921,
			-2041880 when 2922,
			-2042611 when 2923,
			-2043338 when 2924,
			-2044059 when 2925,
			-2044776 when 2926,
			-2045488 when 2927,
			-2046196 when 2928,
			-2046898 when 2929,
			-2047596 when 2930,
			-2048289 when 2931,
			-2048977 when 2932,
			-2049660 when 2933,
			-2050338 when 2934,
			-2051012 when 2935,
			-2051680 when 2936,
			-2052344 when 2937,
			-2053003 when 2938,
			-2053657 when 2939,
			-2054307 when 2940,
			-2054951 when 2941,
			-2055591 when 2942,
			-2056226 when 2943,
			-2056856 when 2944,
			-2057481 when 2945,
			-2058101 when 2946,
			-2058717 when 2947,
			-2059327 when 2948,
			-2059933 when 2949,
			-2060534 when 2950,
			-2061130 when 2951,
			-2061722 when 2952,
			-2062308 when 2953,
			-2062890 when 2954,
			-2063466 when 2955,
			-2064038 when 2956,
			-2064605 when 2957,
			-2065167 when 2958,
			-2065725 when 2959,
			-2066277 when 2960,
			-2066825 when 2961,
			-2067367 when 2962,
			-2067905 when 2963,
			-2068438 when 2964,
			-2068966 when 2965,
			-2069489 when 2966,
			-2070008 when 2967,
			-2070521 when 2968,
			-2071030 when 2969,
			-2071533 when 2970,
			-2072032 when 2971,
			-2072526 when 2972,
			-2073015 when 2973,
			-2073500 when 2974,
			-2073979 when 2975,
			-2074453 when 2976,
			-2074923 when 2977,
			-2075388 when 2978,
			-2075848 when 2979,
			-2076303 when 2980,
			-2076753 when 2981,
			-2077198 when 2982,
			-2077638 when 2983,
			-2078073 when 2984,
			-2078504 when 2985,
			-2078930 when 2986,
			-2079350 when 2987,
			-2079766 when 2988,
			-2080177 when 2989,
			-2080583 when 2990,
			-2080984 when 2991,
			-2081380 when 2992,
			-2081772 when 2993,
			-2082158 when 2994,
			-2082540 when 2995,
			-2082916 when 2996,
			-2083288 when 2997,
			-2083655 when 2998,
			-2084017 when 2999,
			-2084374 when 3000,
			-2084726 when 3001,
			-2085073 when 3002,
			-2085416 when 3003,
			-2085753 when 3004,
			-2086086 when 3005,
			-2086413 when 3006,
			-2086736 when 3007,
			-2087054 when 3008,
			-2087367 when 3009,
			-2087674 when 3010,
			-2087977 when 3011,
			-2088276 when 3012,
			-2088569 when 3013,
			-2088857 when 3014,
			-2089141 when 3015,
			-2089419 when 3016,
			-2089693 when 3017,
			-2089961 when 3018,
			-2090225 when 3019,
			-2090484 when 3020,
			-2090738 when 3021,
			-2090987 when 3022,
			-2091231 when 3023,
			-2091470 when 3024,
			-2091704 when 3025,
			-2091933 when 3026,
			-2092157 when 3027,
			-2092377 when 3028,
			-2092591 when 3029,
			-2092801 when 3030,
			-2093006 when 3031,
			-2093205 when 3032,
			-2093400 when 3033,
			-2093590 when 3034,
			-2093775 when 3035,
			-2093955 when 3036,
			-2094130 when 3037,
			-2094300 when 3038,
			-2094466 when 3039,
			-2094626 when 3040,
			-2094781 when 3041,
			-2094932 when 3042,
			-2095077 when 3043,
			-2095218 when 3044,
			-2095354 when 3045,
			-2095484 when 3046,
			-2095610 when 3047,
			-2095731 when 3048,
			-2095847 when 3049,
			-2095958 when 3050,
			-2096064 when 3051,
			-2096165 when 3052,
			-2096261 when 3053,
			-2096353 when 3054,
			-2096439 when 3055,
			-2096520 when 3056,
			-2096597 when 3057,
			-2096668 when 3058,
			-2096735 when 3059,
			-2096797 when 3060,
			-2096853 when 3061,
			-2096905 when 3062,
			-2096952 when 3063,
			-2096994 when 3064,
			-2097031 when 3065,
			-2097063 when 3066,
			-2097090 when 3067,
			-2097113 when 3068,
			-2097130 when 3069,
			-2097142 when 3070,
			-2097150 when 3071,
			-2097152 when 3072,
			-2097150 when 3073,
			-2097142 when 3074,
			-2097130 when 3075,
			-2097113 when 3076,
			-2097090 when 3077,
			-2097063 when 3078,
			-2097031 when 3079,
			-2096994 when 3080,
			-2096952 when 3081,
			-2096905 when 3082,
			-2096853 when 3083,
			-2096797 when 3084,
			-2096735 when 3085,
			-2096668 when 3086,
			-2096597 when 3087,
			-2096520 when 3088,
			-2096439 when 3089,
			-2096353 when 3090,
			-2096261 when 3091,
			-2096165 when 3092,
			-2096064 when 3093,
			-2095958 when 3094,
			-2095847 when 3095,
			-2095731 when 3096,
			-2095610 when 3097,
			-2095484 when 3098,
			-2095354 when 3099,
			-2095218 when 3100,
			-2095077 when 3101,
			-2094932 when 3102,
			-2094781 when 3103,
			-2094626 when 3104,
			-2094466 when 3105,
			-2094300 when 3106,
			-2094130 when 3107,
			-2093955 when 3108,
			-2093775 when 3109,
			-2093590 when 3110,
			-2093400 when 3111,
			-2093205 when 3112,
			-2093006 when 3113,
			-2092801 when 3114,
			-2092591 when 3115,
			-2092377 when 3116,
			-2092157 when 3117,
			-2091933 when 3118,
			-2091704 when 3119,
			-2091470 when 3120,
			-2091231 when 3121,
			-2090987 when 3122,
			-2090738 when 3123,
			-2090484 when 3124,
			-2090225 when 3125,
			-2089961 when 3126,
			-2089693 when 3127,
			-2089419 when 3128,
			-2089141 when 3129,
			-2088857 when 3130,
			-2088569 when 3131,
			-2088276 when 3132,
			-2087977 when 3133,
			-2087674 when 3134,
			-2087367 when 3135,
			-2087054 when 3136,
			-2086736 when 3137,
			-2086413 when 3138,
			-2086086 when 3139,
			-2085753 when 3140,
			-2085416 when 3141,
			-2085073 when 3142,
			-2084726 when 3143,
			-2084374 when 3144,
			-2084017 when 3145,
			-2083655 when 3146,
			-2083288 when 3147,
			-2082916 when 3148,
			-2082540 when 3149,
			-2082158 when 3150,
			-2081772 when 3151,
			-2081380 when 3152,
			-2080984 when 3153,
			-2080583 when 3154,
			-2080177 when 3155,
			-2079766 when 3156,
			-2079350 when 3157,
			-2078930 when 3158,
			-2078504 when 3159,
			-2078073 when 3160,
			-2077638 when 3161,
			-2077198 when 3162,
			-2076753 when 3163,
			-2076303 when 3164,
			-2075848 when 3165,
			-2075388 when 3166,
			-2074923 when 3167,
			-2074453 when 3168,
			-2073979 when 3169,
			-2073500 when 3170,
			-2073015 when 3171,
			-2072526 when 3172,
			-2072032 when 3173,
			-2071533 when 3174,
			-2071030 when 3175,
			-2070521 when 3176,
			-2070008 when 3177,
			-2069489 when 3178,
			-2068966 when 3179,
			-2068438 when 3180,
			-2067905 when 3181,
			-2067367 when 3182,
			-2066825 when 3183,
			-2066277 when 3184,
			-2065725 when 3185,
			-2065167 when 3186,
			-2064605 when 3187,
			-2064038 when 3188,
			-2063466 when 3189,
			-2062890 when 3190,
			-2062308 when 3191,
			-2061722 when 3192,
			-2061130 when 3193,
			-2060534 when 3194,
			-2059933 when 3195,
			-2059327 when 3196,
			-2058717 when 3197,
			-2058101 when 3198,
			-2057481 when 3199,
			-2056856 when 3200,
			-2056226 when 3201,
			-2055591 when 3202,
			-2054951 when 3203,
			-2054307 when 3204,
			-2053657 when 3205,
			-2053003 when 3206,
			-2052344 when 3207,
			-2051680 when 3208,
			-2051012 when 3209,
			-2050338 when 3210,
			-2049660 when 3211,
			-2048977 when 3212,
			-2048289 when 3213,
			-2047596 when 3214,
			-2046898 when 3215,
			-2046196 when 3216,
			-2045488 when 3217,
			-2044776 when 3218,
			-2044059 when 3219,
			-2043338 when 3220,
			-2042611 when 3221,
			-2041880 when 3222,
			-2041144 when 3223,
			-2040403 when 3224,
			-2039657 when 3225,
			-2038907 when 3226,
			-2038151 when 3227,
			-2037391 when 3228,
			-2036626 when 3229,
			-2035857 when 3230,
			-2035082 when 3231,
			-2034303 when 3232,
			-2033519 when 3233,
			-2032730 when 3234,
			-2031936 when 3235,
			-2031138 when 3236,
			-2030335 when 3237,
			-2029527 when 3238,
			-2028714 when 3239,
			-2027897 when 3240,
			-2027074 when 3241,
			-2026247 when 3242,
			-2025415 when 3243,
			-2024579 when 3244,
			-2023738 when 3245,
			-2022891 when 3246,
			-2022041 when 3247,
			-2021185 when 3248,
			-2020325 when 3249,
			-2019459 when 3250,
			-2018589 when 3251,
			-2017715 when 3252,
			-2016835 when 3253,
			-2015951 when 3254,
			-2015062 when 3255,
			-2014169 when 3256,
			-2013270 when 3257,
			-2012367 when 3258,
			-2011459 when 3259,
			-2010547 when 3260,
			-2009630 when 3261,
			-2008708 when 3262,
			-2007781 when 3263,
			-2006849 when 3264,
			-2005913 when 3265,
			-2004972 when 3266,
			-2004027 when 3267,
			-2003076 when 3268,
			-2002121 when 3269,
			-2001161 when 3270,
			-2000197 when 3271,
			-1999228 when 3272,
			-1998254 when 3273,
			-1997275 when 3274,
			-1996292 when 3275,
			-1995304 when 3276,
			-1994311 when 3277,
			-1993314 when 3278,
			-1992312 when 3279,
			-1991305 when 3280,
			-1990293 when 3281,
			-1989277 when 3282,
			-1988257 when 3283,
			-1987231 when 3284,
			-1986201 when 3285,
			-1985166 when 3286,
			-1984126 when 3287,
			-1983082 when 3288,
			-1982033 when 3289,
			-1980980 when 3290,
			-1979922 when 3291,
			-1978859 when 3292,
			-1977791 when 3293,
			-1976719 when 3294,
			-1975642 when 3295,
			-1974561 when 3296,
			-1973475 when 3297,
			-1972384 when 3298,
			-1971289 when 3299,
			-1970189 when 3300,
			-1969084 when 3301,
			-1967975 when 3302,
			-1966861 when 3303,
			-1965742 when 3304,
			-1964619 when 3305,
			-1963491 when 3306,
			-1962359 when 3307,
			-1961222 when 3308,
			-1960080 when 3309,
			-1958934 when 3310,
			-1957783 when 3311,
			-1956628 when 3312,
			-1955468 when 3313,
			-1954303 when 3314,
			-1953134 when 3315,
			-1951960 when 3316,
			-1950781 when 3317,
			-1949598 when 3318,
			-1948411 when 3319,
			-1947218 when 3320,
			-1946022 when 3321,
			-1944820 when 3322,
			-1943614 when 3323,
			-1942404 when 3324,
			-1941189 when 3325,
			-1939969 when 3326,
			-1938745 when 3327,
			-1937516 when 3328,
			-1936282 when 3329,
			-1935045 when 3330,
			-1933802 when 3331,
			-1932555 when 3332,
			-1931303 when 3333,
			-1930047 when 3334,
			-1928787 when 3335,
			-1927521 when 3336,
			-1926252 when 3337,
			-1924977 when 3338,
			-1923699 when 3339,
			-1922415 when 3340,
			-1921127 when 3341,
			-1919835 when 3342,
			-1918538 when 3343,
			-1917237 when 3344,
			-1915931 when 3345,
			-1914620 when 3346,
			-1913306 when 3347,
			-1911986 when 3348,
			-1910662 when 3349,
			-1909334 when 3350,
			-1908001 when 3351,
			-1906663 when 3352,
			-1905322 when 3353,
			-1903975 when 3354,
			-1902624 when 3355,
			-1901269 when 3356,
			-1899909 when 3357,
			-1898545 when 3358,
			-1897176 when 3359,
			-1895803 when 3360,
			-1894425 when 3361,
			-1893043 when 3362,
			-1891657 when 3363,
			-1890266 when 3364,
			-1888870 when 3365,
			-1887470 when 3366,
			-1886066 when 3367,
			-1884657 when 3368,
			-1883244 when 3369,
			-1881826 when 3370,
			-1880404 when 3371,
			-1878977 when 3372,
			-1877546 when 3373,
			-1876111 when 3374,
			-1874671 when 3375,
			-1873227 when 3376,
			-1871779 when 3377,
			-1870326 when 3378,
			-1868868 when 3379,
			-1867406 when 3380,
			-1865940 when 3381,
			-1864470 when 3382,
			-1862995 when 3383,
			-1861515 when 3384,
			-1860031 when 3385,
			-1858543 when 3386,
			-1857051 when 3387,
			-1855554 when 3388,
			-1854053 when 3389,
			-1852547 when 3390,
			-1851037 when 3391,
			-1849523 when 3392,
			-1848004 when 3393,
			-1846481 when 3394,
			-1844954 when 3395,
			-1843422 when 3396,
			-1841886 when 3397,
			-1840346 when 3398,
			-1838801 when 3399,
			-1837252 when 3400,
			-1835699 when 3401,
			-1834141 when 3402,
			-1832579 when 3403,
			-1831013 when 3404,
			-1829442 when 3405,
			-1827867 when 3406,
			-1826288 when 3407,
			-1824705 when 3408,
			-1823117 when 3409,
			-1821525 when 3410,
			-1819928 when 3411,
			-1818328 when 3412,
			-1816723 when 3413,
			-1815114 when 3414,
			-1813500 when 3415,
			-1811882 when 3416,
			-1810260 when 3417,
			-1808634 when 3418,
			-1807004 when 3419,
			-1805369 when 3420,
			-1803730 when 3421,
			-1802087 when 3422,
			-1800439 when 3423,
			-1798787 when 3424,
			-1797131 when 3425,
			-1795471 when 3426,
			-1793807 when 3427,
			-1792138 when 3428,
			-1790465 when 3429,
			-1788788 when 3430,
			-1787107 when 3431,
			-1785421 when 3432,
			-1783732 when 3433,
			-1782038 when 3434,
			-1780340 when 3435,
			-1778637 when 3436,
			-1776931 when 3437,
			-1775220 when 3438,
			-1773505 when 3439,
			-1771786 when 3440,
			-1770063 when 3441,
			-1768336 when 3442,
			-1766604 when 3443,
			-1764869 when 3444,
			-1763129 when 3445,
			-1761385 when 3446,
			-1759637 when 3447,
			-1757885 when 3448,
			-1756128 when 3449,
			-1754368 when 3450,
			-1752603 when 3451,
			-1750834 when 3452,
			-1749061 when 3453,
			-1747284 when 3454,
			-1745503 when 3455,
			-1743718 when 3456,
			-1741929 when 3457,
			-1740135 when 3458,
			-1738338 when 3459,
			-1736536 when 3460,
			-1734731 when 3461,
			-1732921 when 3462,
			-1731107 when 3463,
			-1729289 when 3464,
			-1727467 when 3465,
			-1725641 when 3466,
			-1723811 when 3467,
			-1721977 when 3468,
			-1720139 when 3469,
			-1718296 when 3470,
			-1716450 when 3471,
			-1714600 when 3472,
			-1712745 when 3473,
			-1710887 when 3474,
			-1709024 when 3475,
			-1707158 when 3476,
			-1705287 when 3477,
			-1703413 when 3478,
			-1701534 when 3479,
			-1699652 when 3480,
			-1697765 when 3481,
			-1695875 when 3482,
			-1693980 when 3483,
			-1692082 when 3484,
			-1690180 when 3485,
			-1688273 when 3486,
			-1686363 when 3487,
			-1684448 when 3488,
			-1682530 when 3489,
			-1680608 when 3490,
			-1678681 when 3491,
			-1676751 when 3492,
			-1674817 when 3493,
			-1672879 when 3494,
			-1670937 when 3495,
			-1668991 when 3496,
			-1667041 when 3497,
			-1665087 when 3498,
			-1663130 when 3499,
			-1661168 when 3500,
			-1659202 when 3501,
			-1657233 when 3502,
			-1655260 when 3503,
			-1653282 when 3504,
			-1651301 when 3505,
			-1649316 when 3506,
			-1647327 when 3507,
			-1645334 when 3508,
			-1643338 when 3509,
			-1641337 when 3510,
			-1639333 when 3511,
			-1637325 when 3512,
			-1635313 when 3513,
			-1633297 when 3514,
			-1631277 when 3515,
			-1629253 when 3516,
			-1627226 when 3517,
			-1625194 when 3518,
			-1623159 when 3519,
			-1621120 when 3520,
			-1619078 when 3521,
			-1617031 when 3522,
			-1614981 when 3523,
			-1612927 when 3524,
			-1610869 when 3525,
			-1608807 when 3526,
			-1606741 when 3527,
			-1604672 when 3528,
			-1602599 when 3529,
			-1600522 when 3530,
			-1598441 when 3531,
			-1596357 when 3532,
			-1594269 when 3533,
			-1592177 when 3534,
			-1590081 when 3535,
			-1587982 when 3536,
			-1585879 when 3537,
			-1583772 when 3538,
			-1581662 when 3539,
			-1579547 when 3540,
			-1577429 when 3541,
			-1575307 when 3542,
			-1573182 when 3543,
			-1571053 when 3544,
			-1568920 when 3545,
			-1566784 when 3546,
			-1564643 when 3547,
			-1562499 when 3548,
			-1560352 when 3549,
			-1558201 when 3550,
			-1556046 when 3551,
			-1553887 when 3552,
			-1551725 when 3553,
			-1549559 when 3554,
			-1547390 when 3555,
			-1545216 when 3556,
			-1543040 when 3557,
			-1540859 when 3558,
			-1538675 when 3559,
			-1536487 when 3560,
			-1534296 when 3561,
			-1532101 when 3562,
			-1529903 when 3563,
			-1527701 when 3564,
			-1525495 when 3565,
			-1523286 when 3566,
			-1521073 when 3567,
			-1518856 when 3568,
			-1516636 when 3569,
			-1514413 when 3570,
			-1512185 when 3571,
			-1509955 when 3572,
			-1507720 when 3573,
			-1505483 when 3574,
			-1503241 when 3575,
			-1500996 when 3576,
			-1498748 when 3577,
			-1496496 when 3578,
			-1494240 when 3579,
			-1491981 when 3580,
			-1489719 when 3581,
			-1487453 when 3582,
			-1485183 when 3583,
			-1482910 when 3584,
			-1480634 when 3585,
			-1478354 when 3586,
			-1476070 when 3587,
			-1473784 when 3588,
			-1471493 when 3589,
			-1469199 when 3590,
			-1466902 when 3591,
			-1464601 when 3592,
			-1462297 when 3593,
			-1459989 when 3594,
			-1457678 when 3595,
			-1455364 when 3596,
			-1453046 when 3597,
			-1450724 when 3598,
			-1448400 when 3599,
			-1446071 when 3600,
			-1443740 when 3601,
			-1441405 when 3602,
			-1439066 when 3603,
			-1436725 when 3604,
			-1434379 when 3605,
			-1432031 when 3606,
			-1429679 when 3607,
			-1427324 when 3608,
			-1424965 when 3609,
			-1422603 when 3610,
			-1420238 when 3611,
			-1417869 when 3612,
			-1415497 when 3613,
			-1413122 when 3614,
			-1410743 when 3615,
			-1408361 when 3616,
			-1405976 when 3617,
			-1403587 when 3618,
			-1401195 when 3619,
			-1398800 when 3620,
			-1396402 when 3621,
			-1394000 when 3622,
			-1391595 when 3623,
			-1389187 when 3624,
			-1386775 when 3625,
			-1384360 when 3626,
			-1381942 when 3627,
			-1379521 when 3628,
			-1377096 when 3629,
			-1374668 when 3630,
			-1372237 when 3631,
			-1369803 when 3632,
			-1367365 when 3633,
			-1364924 when 3634,
			-1362480 when 3635,
			-1360033 when 3636,
			-1357583 when 3637,
			-1355129 when 3638,
			-1352673 when 3639,
			-1350213 when 3640,
			-1347749 when 3641,
			-1345283 when 3642,
			-1342814 when 3643,
			-1340341 when 3644,
			-1337865 when 3645,
			-1335386 when 3646,
			-1332904 when 3647,
			-1330419 when 3648,
			-1327931 when 3649,
			-1325439 when 3650,
			-1322945 when 3651,
			-1320447 when 3652,
			-1317946 when 3653,
			-1315442 when 3654,
			-1312935 when 3655,
			-1310425 when 3656,
			-1307912 when 3657,
			-1305396 when 3658,
			-1302877 when 3659,
			-1300354 when 3660,
			-1297829 when 3661,
			-1295300 when 3662,
			-1292769 when 3663,
			-1290234 when 3664,
			-1287697 when 3665,
			-1285156 when 3666,
			-1282612 when 3667,
			-1280066 when 3668,
			-1277516 when 3669,
			-1274963 when 3670,
			-1272407 when 3671,
			-1269849 when 3672,
			-1267287 when 3673,
			-1264722 when 3674,
			-1262155 when 3675,
			-1259584 when 3676,
			-1257010 when 3677,
			-1254434 when 3678,
			-1251854 when 3679,
			-1249272 when 3680,
			-1246687 when 3681,
			-1244098 when 3682,
			-1241507 when 3683,
			-1238913 when 3684,
			-1236316 when 3685,
			-1233716 when 3686,
			-1231113 when 3687,
			-1228507 when 3688,
			-1225898 when 3689,
			-1223287 when 3690,
			-1220672 when 3691,
			-1218055 when 3692,
			-1215435 when 3693,
			-1212812 when 3694,
			-1210186 when 3695,
			-1207557 when 3696,
			-1204926 when 3697,
			-1202291 when 3698,
			-1199654 when 3699,
			-1197014 when 3700,
			-1194371 when 3701,
			-1191725 when 3702,
			-1189077 when 3703,
			-1186426 when 3704,
			-1183772 when 3705,
			-1181115 when 3706,
			-1178455 when 3707,
			-1175793 when 3708,
			-1173127 when 3709,
			-1170459 when 3710,
			-1167789 when 3711,
			-1165115 when 3712,
			-1162439 when 3713,
			-1159760 when 3714,
			-1157078 when 3715,
			-1154394 when 3716,
			-1151707 when 3717,
			-1149017 when 3718,
			-1146325 when 3719,
			-1143629 when 3720,
			-1140931 when 3721,
			-1138231 when 3722,
			-1135528 when 3723,
			-1132822 when 3724,
			-1130113 when 3725,
			-1127402 when 3726,
			-1124688 when 3727,
			-1121971 when 3728,
			-1119252 when 3729,
			-1116530 when 3730,
			-1113806 when 3731,
			-1111079 when 3732,
			-1108349 when 3733,
			-1105617 when 3734,
			-1102882 when 3735,
			-1100144 when 3736,
			-1097404 when 3737,
			-1094662 when 3738,
			-1091916 when 3739,
			-1089168 when 3740,
			-1086418 when 3741,
			-1083665 when 3742,
			-1080910 when 3743,
			-1078152 when 3744,
			-1075391 when 3745,
			-1072628 when 3746,
			-1069862 when 3747,
			-1067094 when 3748,
			-1064323 when 3749,
			-1061550 when 3750,
			-1058775 when 3751,
			-1055997 when 3752,
			-1053216 when 3753,
			-1050433 when 3754,
			-1047647 when 3755,
			-1044859 when 3756,
			-1042069 when 3757,
			-1039276 when 3758,
			-1036480 when 3759,
			-1033682 when 3760,
			-1030882 when 3761,
			-1028079 when 3762,
			-1025274 when 3763,
			-1022467 when 3764,
			-1019657 when 3765,
			-1016845 when 3766,
			-1014030 when 3767,
			-1011213 when 3768,
			-1008393 when 3769,
			-1005571 when 3770,
			-1002747 when 3771,
			-999920 when 3772,
			-997092 when 3773,
			-994260 when 3774,
			-991427 when 3775,
			-988591 when 3776,
			-985752 when 3777,
			-982912 when 3778,
			-980069 when 3779,
			-977224 when 3780,
			-974376 when 3781,
			-971526 when 3782,
			-968674 when 3783,
			-965820 when 3784,
			-962963 when 3785,
			-960104 when 3786,
			-957243 when 3787,
			-954379 when 3788,
			-951514 when 3789,
			-948646 when 3790,
			-945776 when 3791,
			-942903 when 3792,
			-940029 when 3793,
			-937152 when 3794,
			-934273 when 3795,
			-931392 when 3796,
			-928508 when 3797,
			-925623 when 3798,
			-922735 when 3799,
			-919845 when 3800,
			-916953 when 3801,
			-914059 when 3802,
			-911162 when 3803,
			-908264 when 3804,
			-905363 when 3805,
			-902460 when 3806,
			-899555 when 3807,
			-896648 when 3808,
			-893739 when 3809,
			-890828 when 3810,
			-887914 when 3811,
			-884999 when 3812,
			-882081 when 3813,
			-879162 when 3814,
			-876240 when 3815,
			-873316 when 3816,
			-870390 when 3817,
			-867462 when 3818,
			-864533 when 3819,
			-861601 when 3820,
			-858667 when 3821,
			-855731 when 3822,
			-852793 when 3823,
			-849853 when 3824,
			-846911 when 3825,
			-843967 when 3826,
			-841021 when 3827,
			-838073 when 3828,
			-835123 when 3829,
			-832171 when 3830,
			-829217 when 3831,
			-826261 when 3832,
			-823303 when 3833,
			-820344 when 3834,
			-817382 when 3835,
			-814419 when 3836,
			-811453 when 3837,
			-808486 when 3838,
			-805516 when 3839,
			-802545 when 3840,
			-799572 when 3841,
			-796597 when 3842,
			-793621 when 3843,
			-790642 when 3844,
			-787661 when 3845,
			-784679 when 3846,
			-781695 when 3847,
			-778709 when 3848,
			-775721 when 3849,
			-772731 when 3850,
			-769739 when 3851,
			-766746 when 3852,
			-763751 when 3853,
			-760754 when 3854,
			-757755 when 3855,
			-754755 when 3856,
			-751752 when 3857,
			-748748 when 3858,
			-745742 when 3859,
			-742735 when 3860,
			-739725 when 3861,
			-736714 when 3862,
			-733701 when 3863,
			-730687 when 3864,
			-727671 when 3865,
			-724653 when 3866,
			-721633 when 3867,
			-718612 when 3868,
			-715589 when 3869,
			-712564 when 3870,
			-709537 when 3871,
			-706509 when 3872,
			-703479 when 3873,
			-700448 when 3874,
			-697415 when 3875,
			-694380 when 3876,
			-691344 when 3877,
			-688306 when 3878,
			-685266 when 3879,
			-682225 when 3880,
			-679182 when 3881,
			-676138 when 3882,
			-673092 when 3883,
			-670044 when 3884,
			-666995 when 3885,
			-663944 when 3886,
			-660892 when 3887,
			-657838 when 3888,
			-654783 when 3889,
			-651726 when 3890,
			-648667 when 3891,
			-645607 when 3892,
			-642546 when 3893,
			-639483 when 3894,
			-636418 when 3895,
			-633352 when 3896,
			-630285 when 3897,
			-627216 when 3898,
			-624145 when 3899,
			-621073 when 3900,
			-618000 when 3901,
			-614925 when 3902,
			-611849 when 3903,
			-608771 when 3904,
			-605692 when 3905,
			-602611 when 3906,
			-599529 when 3907,
			-596446 when 3908,
			-593361 when 3909,
			-590275 when 3910,
			-587187 when 3911,
			-584098 when 3912,
			-581008 when 3913,
			-577916 when 3914,
			-574823 when 3915,
			-571728 when 3916,
			-568633 when 3917,
			-565535 when 3918,
			-562437 when 3919,
			-559337 when 3920,
			-556236 when 3921,
			-553134 when 3922,
			-550030 when 3923,
			-546925 when 3924,
			-543819 when 3925,
			-540711 when 3926,
			-537602 when 3927,
			-534492 when 3928,
			-531381 when 3929,
			-528268 when 3930,
			-525154 when 3931,
			-522039 when 3932,
			-518923 when 3933,
			-515805 when 3934,
			-512686 when 3935,
			-509566 when 3936,
			-506445 when 3937,
			-503323 when 3938,
			-500199 when 3939,
			-497075 when 3940,
			-493949 when 3941,
			-490822 when 3942,
			-487693 when 3943,
			-484564 when 3944,
			-481433 when 3945,
			-478302 when 3946,
			-475169 when 3947,
			-472035 when 3948,
			-468900 when 3949,
			-465764 when 3950,
			-462627 when 3951,
			-459489 when 3952,
			-456349 when 3953,
			-453209 when 3954,
			-450067 when 3955,
			-446925 when 3956,
			-443781 when 3957,
			-440636 when 3958,
			-437491 when 3959,
			-434344 when 3960,
			-431196 when 3961,
			-428048 when 3962,
			-424898 when 3963,
			-421747 when 3964,
			-418595 when 3965,
			-415442 when 3966,
			-412289 when 3967,
			-409134 when 3968,
			-405978 when 3969,
			-402822 when 3970,
			-399664 when 3971,
			-396506 when 3972,
			-393346 when 3973,
			-390186 when 3974,
			-387025 when 3975,
			-383862 when 3976,
			-380699 when 3977,
			-377535 when 3978,
			-374371 when 3979,
			-371205 when 3980,
			-368038 when 3981,
			-364871 when 3982,
			-361702 when 3983,
			-358533 when 3984,
			-355363 when 3985,
			-352192 when 3986,
			-349020 when 3987,
			-345848 when 3988,
			-342675 when 3989,
			-339500 when 3990,
			-336325 when 3991,
			-333150 when 3992,
			-329973 when 3993,
			-326796 when 3994,
			-323618 when 3995,
			-320439 when 3996,
			-317259 when 3997,
			-314079 when 3998,
			-310898 when 3999,
			-307716 when 4000,
			-304534 when 4001,
			-301350 when 4002,
			-298166 when 4003,
			-294982 when 4004,
			-291796 when 4005,
			-288610 when 4006,
			-285424 when 4007,
			-282236 when 4008,
			-279048 when 4009,
			-275859 when 4010,
			-272670 when 4011,
			-269480 when 4012,
			-266289 when 4013,
			-263098 when 4014,
			-259906 when 4015,
			-256714 when 4016,
			-253521 when 4017,
			-250327 when 4018,
			-247133 when 4019,
			-243938 when 4020,
			-240742 when 4021,
			-237546 when 4022,
			-234350 when 4023,
			-231153 when 4024,
			-227955 when 4025,
			-224757 when 4026,
			-221558 when 4027,
			-218359 when 4028,
			-215159 when 4029,
			-211959 when 4030,
			-208758 when 4031,
			-205557 when 4032,
			-202355 when 4033,
			-199153 when 4034,
			-195950 when 4035,
			-192747 when 4036,
			-189543 when 4037,
			-186339 when 4038,
			-183135 when 4039,
			-179930 when 4040,
			-176725 when 4041,
			-173519 when 4042,
			-170313 when 4043,
			-167106 when 4044,
			-163899 when 4045,
			-160692 when 4046,
			-157484 when 4047,
			-154276 when 4048,
			-151068 when 4049,
			-147859 when 4050,
			-144650 when 4051,
			-141440 when 4052,
			-138230 when 4053,
			-135020 when 4054,
			-131810 when 4055,
			-128599 when 4056,
			-125388 when 4057,
			-122176 when 4058,
			-118965 when 4059,
			-115753 when 4060,
			-112541 when 4061,
			-109328 when 4062,
			-106115 when 4063,
			-102902 when 4064,
			-99689 when 4065,
			-96476 when 4066,
			-93262 when 4067,
			-90048 when 4068,
			-86834 when 4069,
			-83620 when 4070,
			-80405 when 4071,
			-77190 when 4072,
			-73975 when 4073,
			-70760 when 4074,
			-67545 when 4075,
			-64330 when 4076,
			-61114 when 4077,
			-57898 when 4078,
			-54683 when 4079,
			-51467 when 4080,
			-48251 when 4081,
			-45034 when 4082,
			-41818 when 4083,
			-38602 when 4084,
			-35385 when 4085,
			-32169 when 4086,
			-28952 when 4087,
			-25735 when 4088,
			-22519 when 4089,
			-19302 when 4090,
			-16085 when 4091,
			-12868 when 4092,
			-9651 when 4093,
			-6434 when 4094,
			-3217 when 4095,
			0 when others;

end rtl;